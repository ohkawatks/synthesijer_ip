library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity AXIHP_AFTRANS is
  port (
    clk : in std_logic;
    reset : in std_logic;
    class_s0_0000_axi_reader_ARADDR_exp : in std_logic_vector(32-1 downto 0);
    class_s0_0000_axi_reader_ARVALID_exp : in std_logic;
    class_s0_0000_axi_reader_ARREADY_exp : out std_logic;
    class_s0_0000_axi_reader_RDATA_exp : out std_logic_vector(32-1 downto 0);
    class_s0_0000_axi_reader_RRESP_exp : out std_logic_vector(2-1 downto 0);
    class_s0_0000_axi_reader_RVALID_exp : out std_logic;
    class_s0_0000_axi_reader_RREADY_exp : in std_logic;
    class_s0_0000_axi_writer_AWADDR_exp : in std_logic_vector(32-1 downto 0);
    class_s0_0000_axi_writer_AWVALID_exp : in std_logic;
    class_s0_0000_axi_writer_AWREADY_exp : out std_logic;
    class_s0_0000_axi_writer_WDATA_exp : in std_logic_vector(32-1 downto 0);
    class_s0_0000_axi_writer_WVALID_exp : in std_logic;
    class_s0_0000_axi_writer_WREADY_exp : out std_logic;
    class_s0_0000_axi_writer_WSTRB_exp : in std_logic_vector(4-1 downto 0);
    class_s0_0000_axi_writer_BRESP_exp : out std_logic_vector(2-1 downto 0);
    class_s0_0000_axi_writer_BVALID_exp : out std_logic;
    class_s0_0000_axi_writer_BREADY_exp : in std_logic;
    class_m0_0002_class_obj_0000_forbid_exp_exp : in std_logic;
    class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp_exp : out std_logic_vector(32-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp_exp : out std_logic_vector(8-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp_exp : out std_logic;
    class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp_exp : in std_logic;
    class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp_exp : out std_logic_vector(3-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp_exp : out std_logic_vector(2-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp_exp : out std_logic_vector(4-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp_exp : out std_logic_vector(3-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_RDATA_exp_exp : in std_logic_vector(32-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_RRESP_exp_exp : in std_logic_vector(2-1 downto 0);
    class_m0_0002_class_obj_0000_axi_reader_RLAST_exp_exp : in std_logic;
    class_m0_0002_class_obj_0000_axi_reader_RVALID_exp_exp : in std_logic;
    class_m0_0002_class_obj_0000_axi_reader_RREADY_exp_exp : out std_logic;
    class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp_exp : out std_logic_vector(32-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp_exp : out std_logic_vector(8-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp_exp : out std_logic;
    class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp_exp : out std_logic_vector(3-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp_exp : out std_logic_vector(2-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp_exp : out std_logic_vector(4-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp_exp : out std_logic_vector(3-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp_exp : in std_logic;
    class_m0_0002_class_obj_0000_axi_writer_WDATA_exp_exp : out std_logic_vector(32-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_WLAST_exp_exp : out std_logic;
    class_m0_0002_class_obj_0000_axi_writer_WVALID_exp_exp : out std_logic;
    class_m0_0002_class_obj_0000_axi_writer_WREADY_exp_exp : in std_logic;
    class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp_exp : out std_logic_vector(4-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_BRESP_exp_exp : in std_logic_vector(2-1 downto 0);
    class_m0_0002_class_obj_0000_axi_writer_BVALID_exp_exp : in std_logic;
    class_m0_0002_class_obj_0000_axi_writer_BREADY_exp_exp : out std_logic
  );
end AXIHP_AFTRANS;

architecture RTL of AXIHP_AFTRANS is

  attribute mark_debug : string;
  attribute keep : string;

  component axi_lite_slave_32
    port (
      clk : in std_logic;
      reset : in std_logic;
      data_length : out std_logic_vector(32-1 downto 0);
      data_address : in std_logic_vector(32-1 downto 0);
      data_din : in std_logic_vector(32-1 downto 0);
      data_dout : out std_logic_vector(32-1 downto 0);
      data_we : in std_logic;
      data_oe : in std_logic;
      axi_reader_ARADDR : in std_logic_vector(32-1 downto 0);
      axi_reader_ARVALID : in std_logic;
      axi_reader_ARREADY : out std_logic;
      axi_reader_RDATA : out std_logic_vector(32-1 downto 0);
      axi_reader_RRESP : out std_logic_vector(2-1 downto 0);
      axi_reader_RVALID : out std_logic;
      axi_reader_RREADY : in std_logic;
      axi_writer_AWADDR : in std_logic_vector(32-1 downto 0);
      axi_writer_AWVALID : in std_logic;
      axi_writer_AWREADY : out std_logic;
      axi_writer_WDATA : in std_logic_vector(32-1 downto 0);
      axi_writer_WVALID : in std_logic;
      axi_writer_WREADY : out std_logic;
      axi_writer_WSTRB : in std_logic_vector(4-1 downto 0);
      axi_writer_BRESP : out std_logic_vector(2-1 downto 0);
      axi_writer_BVALID : out std_logic;
      axi_writer_BREADY : in std_logic
    );
  end component axi_lite_slave_32;
  component synthesijer_lib_axi_AXIMemIface32RTLTest
    port (
      clk : in std_logic;
      reset : in std_logic;
      class_obj_0000_forbid_exp : in std_logic;
      class_obj_0000_axi_reader_ARADDR_exp : out std_logic_vector(32-1 downto 0);
      class_obj_0000_axi_reader_ARLEN_exp : out std_logic_vector(8-1 downto 0);
      class_obj_0000_axi_reader_ARVALID_exp : out std_logic;
      class_obj_0000_axi_reader_ARREADY_exp : in std_logic;
      class_obj_0000_axi_reader_ARSIZE_exp : out std_logic_vector(3-1 downto 0);
      class_obj_0000_axi_reader_ARBURST_exp : out std_logic_vector(2-1 downto 0);
      class_obj_0000_axi_reader_ARCACHE_exp : out std_logic_vector(4-1 downto 0);
      class_obj_0000_axi_reader_ARPROT_exp : out std_logic_vector(3-1 downto 0);
      class_obj_0000_axi_reader_RDATA_exp : in std_logic_vector(32-1 downto 0);
      class_obj_0000_axi_reader_RRESP_exp : in std_logic_vector(2-1 downto 0);
      class_obj_0000_axi_reader_RLAST_exp : in std_logic;
      class_obj_0000_axi_reader_RVALID_exp : in std_logic;
      class_obj_0000_axi_reader_RREADY_exp : out std_logic;
      class_obj_0000_axi_writer_AWADDR_exp : out std_logic_vector(32-1 downto 0);
      class_obj_0000_axi_writer_AWLEN_exp : out std_logic_vector(8-1 downto 0);
      class_obj_0000_axi_writer_AWVALID_exp : out std_logic;
      class_obj_0000_axi_writer_AWSIZE_exp : out std_logic_vector(3-1 downto 0);
      class_obj_0000_axi_writer_AWBURST_exp : out std_logic_vector(2-1 downto 0);
      class_obj_0000_axi_writer_AWCACHE_exp : out std_logic_vector(4-1 downto 0);
      class_obj_0000_axi_writer_AWPROT_exp : out std_logic_vector(3-1 downto 0);
      class_obj_0000_axi_writer_AWREADY_exp : in std_logic;
      class_obj_0000_axi_writer_WDATA_exp : out std_logic_vector(32-1 downto 0);
      class_obj_0000_axi_writer_WLAST_exp : out std_logic;
      class_obj_0000_axi_writer_WVALID_exp : out std_logic;
      class_obj_0000_axi_writer_WREADY_exp : in std_logic;
      class_obj_0000_axi_writer_WSTRB_exp : out std_logic_vector(4-1 downto 0);
      class_obj_0000_axi_writer_BRESP_exp : in std_logic_vector(2-1 downto 0);
      class_obj_0000_axi_writer_BVALID_exp : in std_logic;
      class_obj_0000_axi_writer_BREADY_exp : out std_logic;
      flush_addr : in signed(32-1 downto 0);
      flush_burst : in signed(32-1 downto 0);
      fetch_addr : in signed(32-1 downto 0);
      fetch_burst : in signed(32-1 downto 0);
      read_offset : in signed(32-1 downto 0);
      write_offset : in signed(32-1 downto 0);
      write_data : in signed(32-1 downto 0);
      flush_busy : out std_logic;
      flush_req : in std_logic;
      fetch_busy : out std_logic;
      fetch_req : in std_logic;
      read_return : out signed(32-1 downto 0);
      read_busy : out std_logic;
      read_req : in std_logic;
      write_busy : out std_logic;
      write_req : in std_logic
    );
  end component synthesijer_lib_axi_AXIMemIface32RTLTest;
  component AffineTransform
    port (
      clk : in std_logic;
      reset : in std_logic;
      width_in : in signed(32-1 downto 0);
      width_we : in std_logic;
      width_out : out signed(32-1 downto 0);
      height_in : in signed(32-1 downto 0);
      height_we : in std_logic;
      height_out : out signed(32-1 downto 0);
      inData_address : in signed(32-1 downto 0);
      inData_we : in std_logic;
      inData_oe : in std_logic;
      inData_din : in signed(32-1 downto 0);
      inData_dout : out signed(32-1 downto 0);
      inData_length : out signed(32-1 downto 0);
      outData_address : in signed(32-1 downto 0);
      outData_we : in std_logic;
      outData_oe : in std_logic;
      outData_din : in signed(32-1 downto 0);
      outData_dout : out signed(32-1 downto 0);
      outData_length : out signed(32-1 downto 0);
      cmpData_address : in signed(32-1 downto 0);
      cmpData_we : in std_logic;
      cmpData_oe : in std_logic;
      cmpData_din : in signed(32-1 downto 0);
      cmpData_dout : out signed(32-1 downto 0);
      cmpData_length : out signed(32-1 downto 0);
      mat00_in : in signed(16-1 downto 0);
      mat00_we : in std_logic;
      mat00_out : out signed(16-1 downto 0);
      mat01_in : in signed(16-1 downto 0);
      mat01_we : in std_logic;
      mat01_out : out signed(16-1 downto 0);
      mat02_in : in signed(16-1 downto 0);
      mat02_we : in std_logic;
      mat02_out : out signed(16-1 downto 0);
      mat10_in : in signed(16-1 downto 0);
      mat10_we : in std_logic;
      mat10_out : out signed(16-1 downto 0);
      mat11_in : in signed(16-1 downto 0);
      mat11_we : in std_logic;
      mat11_out : out signed(16-1 downto 0);
      mat12_in : in signed(16-1 downto 0);
      mat12_we : in std_logic;
      mat12_out : out signed(16-1 downto 0);
      modeInterpolation_in : in std_logic;
      modeInterpolation_we : in std_logic;
      modeInterpolation_out : out std_logic;
      modeCompare_in : in std_logic;
      modeCompare_we : in std_logic;
      modeCompare_out : out std_logic;
      diffCompare_in : in signed(32-1 downto 0);
      diffCompare_we : in std_logic;
      diffCompare_out : out signed(32-1 downto 0);
      clear_busy : out std_logic;
      clear_req : in std_logic;
      proc_busy : out std_logic;
      proc_req : in std_logic
    );
  end component AffineTransform;

  signal clk_sig : std_logic;
  signal reset_sig : std_logic;
  signal class_s0_0000_axi_reader_ARADDR_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_reader_ARVALID_exp_sig : std_logic;
  signal class_s0_0000_axi_reader_ARREADY_exp_sig : std_logic;
  signal class_s0_0000_axi_reader_RDATA_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_reader_RRESP_exp_sig : std_logic_vector(2-1 downto 0);
  signal class_s0_0000_axi_reader_RVALID_exp_sig : std_logic;
  signal class_s0_0000_axi_reader_RREADY_exp_sig : std_logic;
  signal class_s0_0000_axi_writer_AWADDR_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_writer_AWVALID_exp_sig : std_logic;
  signal class_s0_0000_axi_writer_AWREADY_exp_sig : std_logic;
  signal class_s0_0000_axi_writer_WDATA_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_writer_WVALID_exp_sig : std_logic;
  signal class_s0_0000_axi_writer_WREADY_exp_sig : std_logic;
  signal class_s0_0000_axi_writer_WSTRB_exp_sig : std_logic_vector(4-1 downto 0);
  signal class_s0_0000_axi_writer_BRESP_exp_sig : std_logic_vector(2-1 downto 0);
  signal class_s0_0000_axi_writer_BVALID_exp_sig : std_logic;
  signal class_s0_0000_axi_writer_BREADY_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_forbid_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp_exp_sig : std_logic_vector(8-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp_exp_sig : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp_exp_sig : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp_exp_sig : std_logic_vector(4-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp_exp_sig : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_RDATA_exp_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_RRESP_exp_exp_sig : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_RLAST_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_RVALID_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_RREADY_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp_exp_sig : std_logic_vector(8-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp_exp_sig : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp_exp_sig : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp_exp_sig : std_logic_vector(4-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp_exp_sig : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WDATA_exp_exp_sig : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_WLAST_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WVALID_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WREADY_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp_exp_sig : std_logic_vector(4-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_BRESP_exp_exp_sig : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_BVALID_exp_exp_sig : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_BREADY_exp_exp_sig : std_logic;

  signal class_s0_0000_clk : std_logic;
  signal class_s0_0000_reset : std_logic;
  signal class_s0_0000_data_length : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_data_address : std_logic_vector(32-1 downto 0) := (others => '0');
  signal class_s0_0000_data_din : std_logic_vector(32-1 downto 0) := (others => '0');
  signal class_s0_0000_data_dout : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_data_we : std_logic := '0';
  signal class_s0_0000_data_oe : std_logic := '0';
  signal class_s0_0000_axi_reader_ARADDR : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_reader_ARVALID : std_logic;
  signal class_s0_0000_axi_reader_ARREADY : std_logic;
  signal class_s0_0000_axi_reader_RDATA : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_reader_RRESP : std_logic_vector(2-1 downto 0);
  signal class_s0_0000_axi_reader_RVALID : std_logic;
  signal class_s0_0000_axi_reader_RREADY : std_logic;
  signal class_s0_0000_axi_writer_AWADDR : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_writer_AWVALID : std_logic;
  signal class_s0_0000_axi_writer_AWREADY : std_logic;
  signal class_s0_0000_axi_writer_WDATA : std_logic_vector(32-1 downto 0);
  signal class_s0_0000_axi_writer_WVALID : std_logic;
  signal class_s0_0000_axi_writer_WREADY : std_logic;
  signal class_s0_0000_axi_writer_WSTRB : std_logic_vector(4-1 downto 0);
  signal class_s0_0000_axi_writer_BRESP : std_logic_vector(2-1 downto 0);
  signal class_s0_0000_axi_writer_BVALID : std_logic;
  signal class_s0_0000_axi_writer_BREADY : std_logic;
  signal class_m0_0002_clk : std_logic;
  signal class_m0_0002_reset : std_logic;
  signal class_m0_0002_class_obj_0000_forbid_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp : std_logic_vector(8-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp : std_logic_vector(4-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_RDATA_exp : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_RRESP_exp : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_reader_RLAST_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_RVALID_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_reader_RREADY_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp : std_logic_vector(8-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp : std_logic_vector(4-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp : std_logic_vector(3-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WDATA_exp : std_logic_vector(32-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_WLAST_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WVALID_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WREADY_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp : std_logic_vector(4-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_BRESP_exp : std_logic_vector(2-1 downto 0);
  signal class_m0_0002_class_obj_0000_axi_writer_BVALID_exp : std_logic;
  signal class_m0_0002_class_obj_0000_axi_writer_BREADY_exp : std_logic;
  signal class_m0_0002_flush_addr : signed(32-1 downto 0) := (others => '0');
  signal class_m0_0002_flush_burst : signed(32-1 downto 0) := (others => '0');
  signal class_m0_0002_fetch_addr : signed(32-1 downto 0) := (others => '0');
  signal class_m0_0002_fetch_burst : signed(32-1 downto 0) := (others => '0');
  signal class_m0_0002_read_offset : signed(32-1 downto 0) := (others => '0');
  signal class_m0_0002_write_offset : signed(32-1 downto 0) := (others => '0');
  signal class_m0_0002_write_data : signed(32-1 downto 0) := (others => '0');
  signal class_m0_0002_flush_busy : std_logic;
  signal class_m0_0002_flush_req : std_logic := '0';
  signal class_m0_0002_fetch_busy : std_logic;
  signal class_m0_0002_fetch_req : std_logic := '0';
  signal class_m0_0002_read_return : signed(32-1 downto 0);
  signal class_m0_0002_read_busy : std_logic;
  signal class_m0_0002_read_req : std_logic := '0';
  signal class_m0_0002_write_busy : std_logic;
  signal class_m0_0002_write_req : std_logic := '0';
  signal class_at_0004_clk : std_logic;
  signal class_at_0004_reset : std_logic;
  signal class_at_0004_width_in : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_width_we : std_logic := '0';
  signal class_at_0004_width_out : signed(32-1 downto 0);
  signal class_at_0004_height_in : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_height_we : std_logic := '0';
  signal class_at_0004_height_out : signed(32-1 downto 0);
  signal class_at_0004_inData_address : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_inData_we : std_logic := '0';
  signal class_at_0004_inData_oe : std_logic := '0';
  signal class_at_0004_inData_din : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_inData_dout : signed(32-1 downto 0);
  signal class_at_0004_inData_length : signed(32-1 downto 0);
  signal class_at_0004_outData_address : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_outData_we : std_logic := '0';
  signal class_at_0004_outData_oe : std_logic := '0';
  signal class_at_0004_outData_din : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_outData_dout : signed(32-1 downto 0);
  signal class_at_0004_outData_length : signed(32-1 downto 0);
  signal class_at_0004_cmpData_address : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_cmpData_we : std_logic := '0';
  signal class_at_0004_cmpData_oe : std_logic := '0';
  signal class_at_0004_cmpData_din : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_cmpData_dout : signed(32-1 downto 0);
  signal class_at_0004_cmpData_length : signed(32-1 downto 0);
  signal class_at_0004_mat00_in : signed(16-1 downto 0) := (others => '0');
  signal class_at_0004_mat00_we : std_logic := '0';
  signal class_at_0004_mat00_out : signed(16-1 downto 0);
  signal class_at_0004_mat01_in : signed(16-1 downto 0) := (others => '0');
  signal class_at_0004_mat01_we : std_logic := '0';
  signal class_at_0004_mat01_out : signed(16-1 downto 0);
  signal class_at_0004_mat02_in : signed(16-1 downto 0) := (others => '0');
  signal class_at_0004_mat02_we : std_logic := '0';
  signal class_at_0004_mat02_out : signed(16-1 downto 0);
  signal class_at_0004_mat10_in : signed(16-1 downto 0) := (others => '0');
  signal class_at_0004_mat10_we : std_logic := '0';
  signal class_at_0004_mat10_out : signed(16-1 downto 0);
  signal class_at_0004_mat11_in : signed(16-1 downto 0) := (others => '0');
  signal class_at_0004_mat11_we : std_logic := '0';
  signal class_at_0004_mat11_out : signed(16-1 downto 0);
  signal class_at_0004_mat12_in : signed(16-1 downto 0) := (others => '0');
  signal class_at_0004_mat12_we : std_logic := '0';
  signal class_at_0004_mat12_out : signed(16-1 downto 0);
  signal class_at_0004_modeInterpolation_in : std_logic := '0';
  signal class_at_0004_modeInterpolation_we : std_logic := '0';
  signal class_at_0004_modeInterpolation_out : std_logic;
  signal class_at_0004_modeCompare_in : std_logic := '0';
  signal class_at_0004_modeCompare_we : std_logic := '0';
  signal class_at_0004_modeCompare_out : std_logic;
  signal class_at_0004_diffCompare_in : signed(32-1 downto 0) := (others => '0');
  signal class_at_0004_diffCompare_we : std_logic := '0';
  signal class_at_0004_diffCompare_out : signed(32-1 downto 0);
  signal class_at_0004_clear_busy : std_logic;
  signal class_at_0004_clear_req : std_logic := '0';
  signal class_at_0004_proc_busy : std_logic;
  signal class_at_0004_proc_req : std_logic := '0';
  signal class_BS_0006 : signed(32-1 downto 0) := X"00000100";
  signal class_counter_0007 : signed(32-1 downto 0) := X"00000000";
  signal class_reset_0008 : std_logic := '1';
  signal run_aftrans_proc_width_0009 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00010 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00011 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_proc_height_0012 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00013 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00014 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00015 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00016 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00017 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00018 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00019 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00020 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00021 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00022 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00023 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00024 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00025 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00026 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00027 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00028 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00029 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00030 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00031 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00032 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00033 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00034 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00035 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00036 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00037 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00038 : signed(16-1 downto 0) := (others => '0');
  signal field_access_00039 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00040 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_src_addr_0042 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00043 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00044 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_size_0045 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00046 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00047 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_offset_0048 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00049 : std_logic := '0';
  signal binary_expr_00063 : std_logic := '0';
  signal binary_expr_00065 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00066 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00051 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00052 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00061 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00062 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_i_0053 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00054 : std_logic := '0';
  signal unary_expr_00055 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_d_0056 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00057 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00058 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00059 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00060 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_i_0067 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00068 : std_logic := '0';
  signal unary_expr_00069 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_d_0070 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00071 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00072 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00073 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00074 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_src_addr_0075 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00076 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00077 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_size_0078 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00079 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00080 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_offset_0081 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00082 : std_logic := '0';
  signal binary_expr_00096 : std_logic := '0';
  signal binary_expr_00098 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00099 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00084 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00085 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00094 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00095 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_i_0086 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00087 : std_logic := '0';
  signal unary_expr_00088 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_d_0089 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00090 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00091 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00092 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00093 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_i_0100 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00101 : std_logic := '0';
  signal unary_expr_00102 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_d_0103 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00104 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00105 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00106 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00107 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_dst_addr_0108 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00109 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00110 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_size_0111 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00112 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00113 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_offset_0114 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00115 : std_logic := '0';
  signal binary_expr_00129 : std_logic := '0';
  signal binary_expr_00139 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00140 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00125 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00126 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00127 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00128 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_i_0116 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00117 : std_logic := '0';
  signal unary_expr_00118 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_d_0119 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00120 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00121 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00122 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_i_0130 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00131 : std_logic := '0';
  signal unary_expr_00132 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_d_0133 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00134 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00135 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00136 : signed(32-1 downto 0) := (others => '0');
  signal run_memcpy_src_addr_0141 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00142 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00143 : signed(32-1 downto 0) := (others => '0');
  signal run_memcpy_dest_addr_0144 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00145 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00146 : signed(32-1 downto 0) := (others => '0');
  signal run_memcpy_size_0147 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00148 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00149 : signed(32-1 downto 0) := (others => '0');
  signal run_memcpy_offset_0150 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00151 : std_logic := '0';
  signal binary_expr_00160 : std_logic := '0';
  signal binary_expr_00162 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00163 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00165 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00166 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00153 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00154 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00156 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00157 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00158 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00159 : signed(32-1 downto 0) := (others => '0');
  signal unary_expr_00167 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00168 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00169 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00170 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00171 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00172 : std_logic := '0';
  signal main_cmd_0173 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00174 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00175 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00198 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00199 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00200 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00201 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00177 : std_logic := '0';
  signal field_access_00178 : std_logic := '0';
  signal field_access_00180 : std_logic := '0';
  signal field_access_00181 : std_logic := '0';
  signal field_access_00183 : std_logic := '0';
  signal field_access_00184 : std_logic := '0';
  signal field_access_00186 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00187 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00188 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00189 : std_logic := '0';
  signal field_access_00190 : std_logic := '0';
  signal field_access_00192 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00193 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00194 : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_proc_busy : std_logic := '0';
  signal run_aftrans_proc_req_flag : std_logic;
  signal run_aftrans_proc_req_local : std_logic := '0';
  signal run_aftrans_Src2In_busy : std_logic := '0';
  signal run_aftrans_Src2In_req_flag : std_logic;
  signal run_aftrans_Src2In_req_local : std_logic := '0';
  signal run_aftrans_Src2Cmp_busy : std_logic := '0';
  signal run_aftrans_Src2Cmp_req_flag : std_logic;
  signal run_aftrans_Src2Cmp_req_local : std_logic := '0';
  signal run_aftrans_Out2Dst_busy : std_logic := '0';
  signal run_aftrans_Out2Dst_req_flag : std_logic;
  signal run_aftrans_Out2Dst_req_local : std_logic := '0';
  signal run_memcpy_busy : std_logic := '0';
  signal run_memcpy_req_flag : std_logic;
  signal run_memcpy_req_local : std_logic := '0';
  type Type_run_aftrans_proc_method is (
    run_aftrans_proc_method_IDLE,
    run_aftrans_proc_method_S_0000,
    run_aftrans_proc_method_S_0001,
    run_aftrans_proc_method_S_0002,
    run_aftrans_proc_method_S_0003,
    run_aftrans_proc_method_S_0004,
    run_aftrans_proc_method_S_0005,
    run_aftrans_proc_method_S_0006,
    run_aftrans_proc_method_S_0007,
    run_aftrans_proc_method_S_0008,
    run_aftrans_proc_method_S_0009,
    run_aftrans_proc_method_S_0010,
    run_aftrans_proc_method_S_0011,
    run_aftrans_proc_method_S_0012,
    run_aftrans_proc_method_S_0013,
    run_aftrans_proc_method_S_0014,
    run_aftrans_proc_method_S_0015,
    run_aftrans_proc_method_S_0016,
    run_aftrans_proc_method_S_0017,
    run_aftrans_proc_method_S_0018,
    run_aftrans_proc_method_S_0019,
    run_aftrans_proc_method_S_0020,
    run_aftrans_proc_method_S_0021,
    run_aftrans_proc_method_S_0022,
    run_aftrans_proc_method_S_0023,
    run_aftrans_proc_method_S_0024,
    run_aftrans_proc_method_S_0025,
    run_aftrans_proc_method_S_0026,
    run_aftrans_proc_method_S_0027,
    run_aftrans_proc_method_S_0028,
    run_aftrans_proc_method_S_0029,
    run_aftrans_proc_method_S_0030,
    run_aftrans_proc_method_S_0031,
    run_aftrans_proc_method_S_0032,
    run_aftrans_proc_method_S_0033,
    run_aftrans_proc_method_S_0034,
    run_aftrans_proc_method_S_0035,
    run_aftrans_proc_method_S_0036,
    run_aftrans_proc_method_S_0037,
    run_aftrans_proc_method_S_0038,
    run_aftrans_proc_method_S_0039,
    run_aftrans_proc_method_S_0040,
    run_aftrans_proc_method_S_0041,
    run_aftrans_proc_method_S_0042,
    run_aftrans_proc_method_S_0043,
    run_aftrans_proc_method_S_0042_body,
    run_aftrans_proc_method_S_0042_wait  
  );
  signal run_aftrans_proc_method : Type_run_aftrans_proc_method := run_aftrans_proc_method_IDLE;
  signal run_aftrans_proc_method_delay : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_proc_req_flag_d : std_logic := '0';
  signal run_aftrans_proc_req_flag_edge : std_logic;
  signal tmp_0001 : std_logic;
  signal tmp_0002 : std_logic;
  signal tmp_0003 : std_logic;
  signal tmp_0004 : std_logic;
  signal proc_ext_call_flag_0042 : std_logic;
  signal tmp_0005 : std_logic;
  signal tmp_0006 : std_logic;
  signal tmp_0007 : std_logic;
  signal tmp_0008 : std_logic;
  signal tmp_0009 : std_logic;
  signal tmp_0010 : std_logic;
  signal tmp_0011 : std_logic;
  signal tmp_0012 : std_logic;
  signal tmp_0013 : signed(16-1 downto 0);
  signal tmp_0014 : signed(16-1 downto 0);
  signal tmp_0015 : signed(16-1 downto 0);
  signal tmp_0016 : signed(16-1 downto 0);
  signal tmp_0017 : signed(16-1 downto 0);
  signal tmp_0018 : signed(16-1 downto 0);
  type Type_run_aftrans_Src2In_method is (
    run_aftrans_Src2In_method_IDLE,
    run_aftrans_Src2In_method_S_0000,
    run_aftrans_Src2In_method_S_0001,
    run_aftrans_Src2In_method_S_0002,
    run_aftrans_Src2In_method_S_0003,
    run_aftrans_Src2In_method_S_0004,
    run_aftrans_Src2In_method_S_0005,
    run_aftrans_Src2In_method_S_0006,
    run_aftrans_Src2In_method_S_0007,
    run_aftrans_Src2In_method_S_0009,
    run_aftrans_Src2In_method_S_0010,
    run_aftrans_Src2In_method_S_0011,
    run_aftrans_Src2In_method_S_0012,
    run_aftrans_Src2In_method_S_0013,
    run_aftrans_Src2In_method_S_0014,
    run_aftrans_Src2In_method_S_0015,
    run_aftrans_Src2In_method_S_0016,
    run_aftrans_Src2In_method_S_0017,
    run_aftrans_Src2In_method_S_0018,
    run_aftrans_Src2In_method_S_0019,
    run_aftrans_Src2In_method_S_0020,
    run_aftrans_Src2In_method_S_0021,
    run_aftrans_Src2In_method_S_0022,
    run_aftrans_Src2In_method_S_0023,
    run_aftrans_Src2In_method_S_0024,
    run_aftrans_Src2In_method_S_0025,
    run_aftrans_Src2In_method_S_0026,
    run_aftrans_Src2In_method_S_0028,
    run_aftrans_Src2In_method_S_0029,
    run_aftrans_Src2In_method_S_0030,
    run_aftrans_Src2In_method_S_0033,
    run_aftrans_Src2In_method_S_0034,
    run_aftrans_Src2In_method_S_0035,
    run_aftrans_Src2In_method_S_0036,
    run_aftrans_Src2In_method_S_0037,
    run_aftrans_Src2In_method_S_0038,
    run_aftrans_Src2In_method_S_0039,
    run_aftrans_Src2In_method_S_0040,
    run_aftrans_Src2In_method_S_0041,
    run_aftrans_Src2In_method_S_0042,
    run_aftrans_Src2In_method_S_0043,
    run_aftrans_Src2In_method_S_0044,
    run_aftrans_Src2In_method_S_0045,
    run_aftrans_Src2In_method_S_0046,
    run_aftrans_Src2In_method_S_0047,
    run_aftrans_Src2In_method_S_0048,
    run_aftrans_Src2In_method_S_0049,
    run_aftrans_Src2In_method_S_0050,
    run_aftrans_Src2In_method_S_0051,
    run_aftrans_Src2In_method_S_0052,
    run_aftrans_Src2In_method_S_0053,
    run_aftrans_Src2In_method_S_0055,
    run_aftrans_Src2In_method_S_0056,
    run_aftrans_Src2In_method_S_0014_body,
    run_aftrans_Src2In_method_S_0014_wait,
    run_aftrans_Src2In_method_S_0022_body,
    run_aftrans_Src2In_method_S_0022_wait,
    run_aftrans_Src2In_method_S_0041_body,
    run_aftrans_Src2In_method_S_0041_wait,
    run_aftrans_Src2In_method_S_0049_body,
    run_aftrans_Src2In_method_S_0049_wait  
  );
  signal run_aftrans_Src2In_method : Type_run_aftrans_Src2In_method := run_aftrans_Src2In_method_IDLE;
  signal run_aftrans_Src2In_method_delay : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2In_req_flag_d : std_logic := '0';
  signal run_aftrans_Src2In_req_flag_edge : std_logic;
  signal tmp_0019 : std_logic;
  signal tmp_0020 : std_logic;
  signal tmp_0021 : std_logic;
  signal tmp_0022 : std_logic;
  signal tmp_0023 : std_logic;
  signal tmp_0024 : std_logic;
  signal fetch_ext_call_flag_0014 : std_logic;
  signal tmp_0025 : std_logic;
  signal tmp_0026 : std_logic;
  signal tmp_0027 : std_logic;
  signal tmp_0028 : std_logic;
  signal tmp_0029 : std_logic;
  signal tmp_0030 : std_logic;
  signal read_ext_call_flag_0022 : std_logic;
  signal tmp_0031 : std_logic;
  signal tmp_0032 : std_logic;
  signal tmp_0033 : std_logic;
  signal tmp_0034 : std_logic;
  signal tmp_0035 : std_logic;
  signal tmp_0036 : std_logic;
  signal fetch_ext_call_flag_0041 : std_logic;
  signal tmp_0037 : std_logic;
  signal tmp_0038 : std_logic;
  signal tmp_0039 : std_logic;
  signal tmp_0040 : std_logic;
  signal tmp_0041 : std_logic;
  signal tmp_0042 : std_logic;
  signal read_ext_call_flag_0049 : std_logic;
  signal tmp_0043 : std_logic;
  signal tmp_0044 : std_logic;
  signal tmp_0045 : std_logic;
  signal tmp_0046 : std_logic;
  signal tmp_0047 : std_logic;
  signal tmp_0048 : std_logic;
  signal tmp_0049 : std_logic;
  signal tmp_0050 : std_logic;
  signal tmp_0051 : std_logic;
  signal tmp_0052 : signed(32-1 downto 0);
  signal tmp_0053 : signed(32-1 downto 0);
  signal tmp_0054 : std_logic;
  signal tmp_0055 : signed(32-1 downto 0);
  signal tmp_0056 : signed(32-1 downto 0);
  signal tmp_0057 : signed(32-1 downto 0);
  signal tmp_0058 : signed(32-1 downto 0);
  signal tmp_0059 : std_logic;
  signal tmp_0060 : signed(32-1 downto 0);
  signal tmp_0061 : signed(32-1 downto 0);
  signal tmp_0062 : std_logic;
  signal tmp_0063 : signed(32-1 downto 0);
  signal tmp_0064 : signed(32-1 downto 0);
  type Type_run_aftrans_Src2Cmp_method is (
    run_aftrans_Src2Cmp_method_IDLE,
    run_aftrans_Src2Cmp_method_S_0000,
    run_aftrans_Src2Cmp_method_S_0001,
    run_aftrans_Src2Cmp_method_S_0002,
    run_aftrans_Src2Cmp_method_S_0003,
    run_aftrans_Src2Cmp_method_S_0004,
    run_aftrans_Src2Cmp_method_S_0005,
    run_aftrans_Src2Cmp_method_S_0006,
    run_aftrans_Src2Cmp_method_S_0007,
    run_aftrans_Src2Cmp_method_S_0009,
    run_aftrans_Src2Cmp_method_S_0010,
    run_aftrans_Src2Cmp_method_S_0011,
    run_aftrans_Src2Cmp_method_S_0012,
    run_aftrans_Src2Cmp_method_S_0013,
    run_aftrans_Src2Cmp_method_S_0014,
    run_aftrans_Src2Cmp_method_S_0015,
    run_aftrans_Src2Cmp_method_S_0016,
    run_aftrans_Src2Cmp_method_S_0017,
    run_aftrans_Src2Cmp_method_S_0018,
    run_aftrans_Src2Cmp_method_S_0019,
    run_aftrans_Src2Cmp_method_S_0020,
    run_aftrans_Src2Cmp_method_S_0021,
    run_aftrans_Src2Cmp_method_S_0022,
    run_aftrans_Src2Cmp_method_S_0023,
    run_aftrans_Src2Cmp_method_S_0024,
    run_aftrans_Src2Cmp_method_S_0025,
    run_aftrans_Src2Cmp_method_S_0026,
    run_aftrans_Src2Cmp_method_S_0028,
    run_aftrans_Src2Cmp_method_S_0029,
    run_aftrans_Src2Cmp_method_S_0030,
    run_aftrans_Src2Cmp_method_S_0033,
    run_aftrans_Src2Cmp_method_S_0034,
    run_aftrans_Src2Cmp_method_S_0035,
    run_aftrans_Src2Cmp_method_S_0036,
    run_aftrans_Src2Cmp_method_S_0037,
    run_aftrans_Src2Cmp_method_S_0038,
    run_aftrans_Src2Cmp_method_S_0039,
    run_aftrans_Src2Cmp_method_S_0040,
    run_aftrans_Src2Cmp_method_S_0041,
    run_aftrans_Src2Cmp_method_S_0042,
    run_aftrans_Src2Cmp_method_S_0043,
    run_aftrans_Src2Cmp_method_S_0044,
    run_aftrans_Src2Cmp_method_S_0045,
    run_aftrans_Src2Cmp_method_S_0046,
    run_aftrans_Src2Cmp_method_S_0047,
    run_aftrans_Src2Cmp_method_S_0048,
    run_aftrans_Src2Cmp_method_S_0049,
    run_aftrans_Src2Cmp_method_S_0050,
    run_aftrans_Src2Cmp_method_S_0051,
    run_aftrans_Src2Cmp_method_S_0052,
    run_aftrans_Src2Cmp_method_S_0053,
    run_aftrans_Src2Cmp_method_S_0055,
    run_aftrans_Src2Cmp_method_S_0056,
    run_aftrans_Src2Cmp_method_S_0014_body,
    run_aftrans_Src2Cmp_method_S_0014_wait,
    run_aftrans_Src2Cmp_method_S_0022_body,
    run_aftrans_Src2Cmp_method_S_0022_wait,
    run_aftrans_Src2Cmp_method_S_0041_body,
    run_aftrans_Src2Cmp_method_S_0041_wait,
    run_aftrans_Src2Cmp_method_S_0049_body,
    run_aftrans_Src2Cmp_method_S_0049_wait  
  );
  signal run_aftrans_Src2Cmp_method : Type_run_aftrans_Src2Cmp_method := run_aftrans_Src2Cmp_method_IDLE;
  signal run_aftrans_Src2Cmp_method_delay : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Src2Cmp_req_flag_d : std_logic := '0';
  signal run_aftrans_Src2Cmp_req_flag_edge : std_logic;
  signal tmp_0065 : std_logic;
  signal tmp_0066 : std_logic;
  signal tmp_0067 : std_logic;
  signal tmp_0068 : std_logic;
  signal tmp_0069 : std_logic;
  signal tmp_0070 : std_logic;
  signal tmp_0071 : std_logic;
  signal tmp_0072 : std_logic;
  signal tmp_0073 : std_logic;
  signal tmp_0074 : std_logic;
  signal tmp_0075 : std_logic;
  signal tmp_0076 : std_logic;
  signal tmp_0077 : std_logic;
  signal tmp_0078 : std_logic;
  signal tmp_0079 : std_logic;
  signal tmp_0080 : std_logic;
  signal tmp_0081 : std_logic;
  signal tmp_0082 : signed(32-1 downto 0);
  signal tmp_0083 : signed(32-1 downto 0);
  signal tmp_0084 : std_logic;
  signal tmp_0085 : signed(32-1 downto 0);
  signal tmp_0086 : signed(32-1 downto 0);
  signal tmp_0087 : signed(32-1 downto 0);
  signal tmp_0088 : signed(32-1 downto 0);
  signal tmp_0089 : std_logic;
  signal tmp_0090 : signed(32-1 downto 0);
  signal tmp_0091 : signed(32-1 downto 0);
  signal tmp_0092 : std_logic;
  signal tmp_0093 : signed(32-1 downto 0);
  signal tmp_0094 : signed(32-1 downto 0);
  type Type_run_aftrans_Out2Dst_method is (
    run_aftrans_Out2Dst_method_IDLE,
    run_aftrans_Out2Dst_method_S_0000,
    run_aftrans_Out2Dst_method_S_0001,
    run_aftrans_Out2Dst_method_S_0002,
    run_aftrans_Out2Dst_method_S_0003,
    run_aftrans_Out2Dst_method_S_0004,
    run_aftrans_Out2Dst_method_S_0005,
    run_aftrans_Out2Dst_method_S_0006,
    run_aftrans_Out2Dst_method_S_0007,
    run_aftrans_Out2Dst_method_S_0009,
    run_aftrans_Out2Dst_method_S_0010,
    run_aftrans_Out2Dst_method_S_0011,
    run_aftrans_Out2Dst_method_S_0012,
    run_aftrans_Out2Dst_method_S_0013,
    run_aftrans_Out2Dst_method_S_0014,
    run_aftrans_Out2Dst_method_S_0015,
    run_aftrans_Out2Dst_method_S_0016,
    run_aftrans_Out2Dst_method_S_0017,
    run_aftrans_Out2Dst_method_S_0018,
    run_aftrans_Out2Dst_method_S_0019,
    run_aftrans_Out2Dst_method_S_0020,
    run_aftrans_Out2Dst_method_S_0021,
    run_aftrans_Out2Dst_method_S_0022,
    run_aftrans_Out2Dst_method_S_0023,
    run_aftrans_Out2Dst_method_S_0024,
    run_aftrans_Out2Dst_method_S_0025,
    run_aftrans_Out2Dst_method_S_0026,
    run_aftrans_Out2Dst_method_S_0027,
    run_aftrans_Out2Dst_method_S_0028,
    run_aftrans_Out2Dst_method_S_0029,
    run_aftrans_Out2Dst_method_S_0032,
    run_aftrans_Out2Dst_method_S_0033,
    run_aftrans_Out2Dst_method_S_0034,
    run_aftrans_Out2Dst_method_S_0035,
    run_aftrans_Out2Dst_method_S_0036,
    run_aftrans_Out2Dst_method_S_0037,
    run_aftrans_Out2Dst_method_S_0038,
    run_aftrans_Out2Dst_method_S_0039,
    run_aftrans_Out2Dst_method_S_0040,
    run_aftrans_Out2Dst_method_S_0041,
    run_aftrans_Out2Dst_method_S_0042,
    run_aftrans_Out2Dst_method_S_0043,
    run_aftrans_Out2Dst_method_S_0044,
    run_aftrans_Out2Dst_method_S_0045,
    run_aftrans_Out2Dst_method_S_0046,
    run_aftrans_Out2Dst_method_S_0047,
    run_aftrans_Out2Dst_method_S_0048,
    run_aftrans_Out2Dst_method_S_0049,
    run_aftrans_Out2Dst_method_S_0050,
    run_aftrans_Out2Dst_method_S_0051,
    run_aftrans_Out2Dst_method_S_0052,
    run_aftrans_Out2Dst_method_S_0053,
    run_aftrans_Out2Dst_method_S_0054,
    run_aftrans_Out2Dst_method_S_0023_body,
    run_aftrans_Out2Dst_method_S_0023_wait,
    run_aftrans_Out2Dst_method_S_0027_body,
    run_aftrans_Out2Dst_method_S_0027_wait,
    run_aftrans_Out2Dst_method_S_0049_body,
    run_aftrans_Out2Dst_method_S_0049_wait,
    run_aftrans_Out2Dst_method_S_0053_body,
    run_aftrans_Out2Dst_method_S_0053_wait  
  );
  signal run_aftrans_Out2Dst_method : Type_run_aftrans_Out2Dst_method := run_aftrans_Out2Dst_method_IDLE;
  signal run_aftrans_Out2Dst_method_delay : signed(32-1 downto 0) := (others => '0');
  signal run_aftrans_Out2Dst_req_flag_d : std_logic := '0';
  signal run_aftrans_Out2Dst_req_flag_edge : std_logic;
  signal tmp_0095 : std_logic;
  signal tmp_0096 : std_logic;
  signal tmp_0097 : std_logic;
  signal tmp_0098 : std_logic;
  signal tmp_0099 : std_logic;
  signal tmp_0100 : std_logic;
  signal tmp_0101 : std_logic;
  signal tmp_0102 : std_logic;
  signal write_ext_call_flag_0023 : std_logic;
  signal tmp_0103 : std_logic;
  signal tmp_0104 : std_logic;
  signal tmp_0105 : std_logic;
  signal tmp_0106 : std_logic;
  signal flush_ext_call_flag_0027 : std_logic;
  signal tmp_0107 : std_logic;
  signal tmp_0108 : std_logic;
  signal tmp_0109 : std_logic;
  signal tmp_0110 : std_logic;
  signal tmp_0111 : std_logic;
  signal tmp_0112 : std_logic;
  signal tmp_0113 : std_logic;
  signal tmp_0114 : std_logic;
  signal write_ext_call_flag_0049 : std_logic;
  signal tmp_0115 : std_logic;
  signal tmp_0116 : std_logic;
  signal tmp_0117 : std_logic;
  signal tmp_0118 : std_logic;
  signal flush_ext_call_flag_0053 : std_logic;
  signal tmp_0119 : std_logic;
  signal tmp_0120 : std_logic;
  signal tmp_0121 : std_logic;
  signal tmp_0122 : std_logic;
  signal tmp_0123 : std_logic;
  signal tmp_0124 : std_logic;
  signal tmp_0125 : std_logic;
  signal tmp_0126 : std_logic;
  signal tmp_0127 : std_logic;
  signal tmp_0128 : std_logic;
  signal tmp_0129 : signed(32-1 downto 0);
  signal tmp_0130 : signed(32-1 downto 0);
  signal tmp_0131 : signed(32-1 downto 0);
  signal tmp_0132 : signed(32-1 downto 0);
  signal tmp_0133 : signed(32-1 downto 0);
  signal tmp_0134 : signed(32-1 downto 0);
  signal tmp_0135 : std_logic;
  signal tmp_0136 : std_logic;
  signal tmp_0137 : signed(32-1 downto 0);
  signal tmp_0138 : signed(32-1 downto 0);
  signal tmp_0139 : signed(32-1 downto 0);
  signal tmp_0140 : signed(32-1 downto 0);
  type Type_run_memcpy_method is (
    run_memcpy_method_IDLE,
    run_memcpy_method_S_0000,
    run_memcpy_method_S_0001,
    run_memcpy_method_S_0002,
    run_memcpy_method_S_0003,
    run_memcpy_method_S_0004,
    run_memcpy_method_S_0005,
    run_memcpy_method_S_0006,
    run_memcpy_method_S_0007,
    run_memcpy_method_S_0008,
    run_memcpy_method_S_0009,
    run_memcpy_method_S_0010,
    run_memcpy_method_S_0012,
    run_memcpy_method_S_0013,
    run_memcpy_method_S_0014,
    run_memcpy_method_S_0015,
    run_memcpy_method_S_0016,
    run_memcpy_method_S_0017,
    run_memcpy_method_S_0018,
    run_memcpy_method_S_0019,
    run_memcpy_method_S_0020,
    run_memcpy_method_S_0021,
    run_memcpy_method_S_0022,
    run_memcpy_method_S_0025,
    run_memcpy_method_S_0026,
    run_memcpy_method_S_0027,
    run_memcpy_method_S_0028,
    run_memcpy_method_S_0029,
    run_memcpy_method_S_0030,
    run_memcpy_method_S_0031,
    run_memcpy_method_S_0032,
    run_memcpy_method_S_0033,
    run_memcpy_method_S_0034,
    run_memcpy_method_S_0035,
    run_memcpy_method_S_0036,
    run_memcpy_method_S_0037,
    run_memcpy_method_S_0017_body,
    run_memcpy_method_S_0017_wait,
    run_memcpy_method_S_0020_body,
    run_memcpy_method_S_0020_wait,
    run_memcpy_method_S_0033_body,
    run_memcpy_method_S_0033_wait,
    run_memcpy_method_S_0036_body,
    run_memcpy_method_S_0036_wait  
  );
  signal run_memcpy_method : Type_run_memcpy_method := run_memcpy_method_IDLE;
  signal run_memcpy_method_delay : signed(32-1 downto 0) := (others => '0');
  signal run_memcpy_req_flag_d : std_logic := '0';
  signal run_memcpy_req_flag_edge : std_logic;
  signal tmp_0141 : std_logic;
  signal tmp_0142 : std_logic;
  signal tmp_0143 : std_logic;
  signal tmp_0144 : std_logic;
  signal tmp_0145 : std_logic;
  signal tmp_0146 : std_logic;
  signal fetch_ext_call_flag_0017 : std_logic;
  signal tmp_0147 : std_logic;
  signal tmp_0148 : std_logic;
  signal tmp_0149 : std_logic;
  signal tmp_0150 : std_logic;
  signal flush_ext_call_flag_0020 : std_logic;
  signal tmp_0151 : std_logic;
  signal tmp_0152 : std_logic;
  signal tmp_0153 : std_logic;
  signal tmp_0154 : std_logic;
  signal tmp_0155 : std_logic;
  signal tmp_0156 : std_logic;
  signal fetch_ext_call_flag_0033 : std_logic;
  signal tmp_0157 : std_logic;
  signal tmp_0158 : std_logic;
  signal tmp_0159 : std_logic;
  signal tmp_0160 : std_logic;
  signal flush_ext_call_flag_0036 : std_logic;
  signal tmp_0161 : std_logic;
  signal tmp_0162 : std_logic;
  signal tmp_0163 : std_logic;
  signal tmp_0164 : std_logic;
  signal tmp_0165 : std_logic;
  signal tmp_0166 : std_logic;
  signal tmp_0167 : std_logic;
  signal tmp_0168 : std_logic;
  signal tmp_0169 : std_logic;
  signal tmp_0170 : signed(32-1 downto 0);
  signal tmp_0171 : signed(32-1 downto 0);
  signal tmp_0172 : signed(32-1 downto 0);
  signal tmp_0173 : signed(32-1 downto 0);
  signal tmp_0174 : signed(32-1 downto 0);
  signal tmp_0175 : signed(32-1 downto 0);
  signal tmp_0176 : std_logic;
  signal tmp_0177 : signed(32-1 downto 0);
  signal tmp_0178 : signed(32-1 downto 0);
  signal tmp_0179 : signed(32-1 downto 0);
  signal tmp_0180 : signed(32-1 downto 0);
  type Type_clock_method is (
    clock_method_IDLE,
    clock_method_S_0000,
    clock_method_S_0001,
    clock_method_S_0002,
    clock_method_S_0003,
    clock_method_S_0004,
    clock_method_S_0005,
    clock_method_S_0006,
    clock_method_S_0008,
    clock_method_S_0009,
    clock_method_S_0010,
    clock_method_S_0011,
    clock_method_S_0012,
    clock_method_S_0013  
  );
  signal clock_method : Type_clock_method := clock_method_IDLE;
  signal clock_method_delay : signed(32-1 downto 0) := (others => '0');
  signal tmp_0181 : std_logic;
  signal tmp_0182 : std_logic;
  signal tmp_0183 : std_logic;
  signal tmp_0184 : std_logic;
  signal tmp_0185 : signed(32-1 downto 0);
  type Type_main_method is (
    main_method_IDLE,
    main_method_S_0000,
    main_method_S_0001,
    main_method_S_0002,
    main_method_S_0003,
    main_method_S_0005,
    main_method_S_0006,
    main_method_S_0007,
    main_method_S_0008,
    main_method_S_0009,
    main_method_S_0010,
    main_method_S_0011,
    main_method_S_0012,
    main_method_S_0013,
    main_method_S_0015,
    main_method_S_0016,
    main_method_S_0017,
    main_method_S_0018,
    main_method_S_0019,
    main_method_S_0020,
    main_method_S_0021,
    main_method_S_0022,
    main_method_S_0023,
    main_method_S_0024,
    main_method_S_0025,
    main_method_S_0026,
    main_method_S_0027,
    main_method_S_0028,
    main_method_S_0029,
    main_method_S_0030,
    main_method_S_0031,
    main_method_S_0032,
    main_method_S_0033,
    main_method_S_0034,
    main_method_S_0035,
    main_method_S_0036,
    main_method_S_0037,
    main_method_S_0038,
    main_method_S_0039,
    main_method_S_0040,
    main_method_S_0041,
    main_method_S_0042,
    main_method_S_0043,
    main_method_S_0044,
    main_method_S_0045,
    main_method_S_0046,
    main_method_S_0047,
    main_method_S_0048,
    main_method_S_0049,
    main_method_S_0050,
    main_method_S_0051,
    main_method_S_0052,
    main_method_S_0053,
    main_method_S_0054,
    main_method_S_0055,
    main_method_S_0056,
    main_method_S_0057,
    main_method_S_0058,
    main_method_S_0059,
    main_method_S_0060,
    main_method_S_0061,
    main_method_S_0062,
    main_method_S_0063,
    main_method_S_0064,
    main_method_S_0065,
    main_method_S_0066,
    main_method_S_0067,
    main_method_S_0069,
    main_method_S_0070,
    main_method_S_0072,
    main_method_S_0018_body,
    main_method_S_0018_wait,
    main_method_S_0025_body,
    main_method_S_0025_wait,
    main_method_S_0032_body,
    main_method_S_0032_wait,
    main_method_S_0039_body,
    main_method_S_0039_wait,
    main_method_S_0050_body,
    main_method_S_0050_wait,
    main_method_S_0057_body,
    main_method_S_0057_wait,
    main_method_S_0060_body,
    main_method_S_0060_wait,
    main_method_S_0063_body,
    main_method_S_0063_wait  
  );
  signal main_method : Type_main_method := main_method_IDLE;
  signal main_method_delay : signed(32-1 downto 0) := (others => '0');
  signal tmp_0186 : std_logic;
  signal tmp_0187 : std_logic;
  signal tmp_0188 : std_logic;
  signal tmp_0189 : std_logic;
  signal tmp_0190 : std_logic;
  signal tmp_0191 : std_logic;
  signal tmp_0192 : std_logic;
  signal tmp_0193 : std_logic;
  signal tmp_0194 : std_logic;
  signal tmp_0195 : std_logic;
  signal run_memcpy_call_flag_0018 : std_logic;
  signal tmp_0196 : std_logic;
  signal tmp_0197 : std_logic;
  signal tmp_0198 : std_logic;
  signal tmp_0199 : std_logic;
  signal run_aftrans_proc_call_flag_0025 : std_logic;
  signal tmp_0200 : std_logic;
  signal tmp_0201 : std_logic;
  signal tmp_0202 : std_logic;
  signal tmp_0203 : std_logic;
  signal run_aftrans_proc_call_flag_0032 : std_logic;
  signal tmp_0204 : std_logic;
  signal tmp_0205 : std_logic;
  signal tmp_0206 : std_logic;
  signal tmp_0207 : std_logic;
  signal run_aftrans_proc_call_flag_0039 : std_logic;
  signal tmp_0208 : std_logic;
  signal tmp_0209 : std_logic;
  signal tmp_0210 : std_logic;
  signal tmp_0211 : std_logic;
  signal run_aftrans_proc_call_flag_0050 : std_logic;
  signal tmp_0212 : std_logic;
  signal tmp_0213 : std_logic;
  signal tmp_0214 : std_logic;
  signal tmp_0215 : std_logic;
  signal run_aftrans_Out2Dst_call_flag_0057 : std_logic;
  signal tmp_0216 : std_logic;
  signal tmp_0217 : std_logic;
  signal tmp_0218 : std_logic;
  signal tmp_0219 : std_logic;
  signal run_aftrans_Src2Cmp_call_flag_0060 : std_logic;
  signal tmp_0220 : std_logic;
  signal tmp_0221 : std_logic;
  signal tmp_0222 : std_logic;
  signal tmp_0223 : std_logic;
  signal run_aftrans_Src2In_call_flag_0063 : std_logic;
  signal tmp_0224 : std_logic;
  signal tmp_0225 : std_logic;
  signal tmp_0226 : std_logic;
  signal tmp_0227 : std_logic;
  signal tmp_0228 : std_logic;

begin

  clk_sig <= clk;
  reset_sig <= reset;
  class_s0_0000_axi_reader_ARADDR_exp_sig <= class_s0_0000_axi_reader_ARADDR_exp;
  class_s0_0000_axi_reader_ARVALID_exp_sig <= class_s0_0000_axi_reader_ARVALID_exp;
  class_s0_0000_axi_reader_ARREADY_exp <= class_s0_0000_axi_reader_ARREADY_exp_sig;
  class_s0_0000_axi_reader_ARREADY_exp_sig <= class_s0_0000_axi_reader_ARREADY;

  class_s0_0000_axi_reader_RDATA_exp <= class_s0_0000_axi_reader_RDATA_exp_sig;
  class_s0_0000_axi_reader_RDATA_exp_sig <= class_s0_0000_axi_reader_RDATA;

  class_s0_0000_axi_reader_RRESP_exp <= class_s0_0000_axi_reader_RRESP_exp_sig;
  class_s0_0000_axi_reader_RRESP_exp_sig <= class_s0_0000_axi_reader_RRESP;

  class_s0_0000_axi_reader_RVALID_exp <= class_s0_0000_axi_reader_RVALID_exp_sig;
  class_s0_0000_axi_reader_RVALID_exp_sig <= class_s0_0000_axi_reader_RVALID;

  class_s0_0000_axi_reader_RREADY_exp_sig <= class_s0_0000_axi_reader_RREADY_exp;
  class_s0_0000_axi_writer_AWADDR_exp_sig <= class_s0_0000_axi_writer_AWADDR_exp;
  class_s0_0000_axi_writer_AWVALID_exp_sig <= class_s0_0000_axi_writer_AWVALID_exp;
  class_s0_0000_axi_writer_AWREADY_exp <= class_s0_0000_axi_writer_AWREADY_exp_sig;
  class_s0_0000_axi_writer_AWREADY_exp_sig <= class_s0_0000_axi_writer_AWREADY;

  class_s0_0000_axi_writer_WDATA_exp_sig <= class_s0_0000_axi_writer_WDATA_exp;
  class_s0_0000_axi_writer_WVALID_exp_sig <= class_s0_0000_axi_writer_WVALID_exp;
  class_s0_0000_axi_writer_WREADY_exp <= class_s0_0000_axi_writer_WREADY_exp_sig;
  class_s0_0000_axi_writer_WREADY_exp_sig <= class_s0_0000_axi_writer_WREADY;

  class_s0_0000_axi_writer_WSTRB_exp_sig <= class_s0_0000_axi_writer_WSTRB_exp;
  class_s0_0000_axi_writer_BRESP_exp <= class_s0_0000_axi_writer_BRESP_exp_sig;
  class_s0_0000_axi_writer_BRESP_exp_sig <= class_s0_0000_axi_writer_BRESP;

  class_s0_0000_axi_writer_BVALID_exp <= class_s0_0000_axi_writer_BVALID_exp_sig;
  class_s0_0000_axi_writer_BVALID_exp_sig <= class_s0_0000_axi_writer_BVALID;

  class_s0_0000_axi_writer_BREADY_exp_sig <= class_s0_0000_axi_writer_BREADY_exp;
  class_m0_0002_class_obj_0000_forbid_exp_exp_sig <= class_m0_0002_class_obj_0000_forbid_exp_exp;
  class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp;

  class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp;

  class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp;

  class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp_exp;
  class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp;

  class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp;

  class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp;

  class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp;

  class_m0_0002_class_obj_0000_axi_reader_RDATA_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_RDATA_exp_exp;
  class_m0_0002_class_obj_0000_axi_reader_RRESP_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_RRESP_exp_exp;
  class_m0_0002_class_obj_0000_axi_reader_RLAST_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_RLAST_exp_exp;
  class_m0_0002_class_obj_0000_axi_reader_RVALID_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_RVALID_exp_exp;
  class_m0_0002_class_obj_0000_axi_reader_RREADY_exp_exp <= class_m0_0002_class_obj_0000_axi_reader_RREADY_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_reader_RREADY_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_reader_RREADY_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp;

  class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp_exp;
  class_m0_0002_class_obj_0000_axi_writer_WDATA_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_WDATA_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_WDATA_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_WDATA_exp;

  class_m0_0002_class_obj_0000_axi_writer_WLAST_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_WLAST_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_WLAST_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_WLAST_exp;

  class_m0_0002_class_obj_0000_axi_writer_WVALID_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_WVALID_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_WVALID_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_WVALID_exp;

  class_m0_0002_class_obj_0000_axi_writer_WREADY_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_WREADY_exp_exp;
  class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp;

  class_m0_0002_class_obj_0000_axi_writer_BRESP_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_BRESP_exp_exp;
  class_m0_0002_class_obj_0000_axi_writer_BVALID_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_BVALID_exp_exp;
  class_m0_0002_class_obj_0000_axi_writer_BREADY_exp_exp <= class_m0_0002_class_obj_0000_axi_writer_BREADY_exp_exp_sig;
  class_m0_0002_class_obj_0000_axi_writer_BREADY_exp_exp_sig <= class_m0_0002_class_obj_0000_axi_writer_BREADY_exp;


  -- expressions
  tmp_0001 <= not run_aftrans_proc_req_flag_d;
  tmp_0002 <= run_aftrans_proc_req_flag and tmp_0001;
  tmp_0003 <= run_aftrans_proc_req_flag or run_aftrans_proc_req_flag_d;
  tmp_0004 <= run_aftrans_proc_req_flag or run_aftrans_proc_req_flag_d;
  tmp_0005 <= '1' when class_at_0004_proc_busy = '0' else '0';
  tmp_0006 <= '1' when class_at_0004_proc_req = '0' else '0';
  tmp_0007 <= tmp_0005 and tmp_0006;
  tmp_0008 <= '1' when tmp_0007 = '1' else '0';
  tmp_0009 <= '1' when run_aftrans_proc_method /= run_aftrans_proc_method_S_0000 else '0';
  tmp_0010 <= '1' when run_aftrans_proc_method /= run_aftrans_proc_method_S_0001 else '0';
  tmp_0011 <= tmp_0010 and run_aftrans_proc_req_flag_edge;
  tmp_0012 <= tmp_0009 and tmp_0011;
  tmp_0013 <= array_access_00017(32 - 16 - 1 downto 0);
  tmp_0014 <= array_access_00021(32 - 16 - 1 downto 0);
  tmp_0015 <= array_access_00025(32 - 16 - 1 downto 0);
  tmp_0016 <= array_access_00029(32 - 16 - 1 downto 0);
  tmp_0017 <= array_access_00033(32 - 16 - 1 downto 0);
  tmp_0018 <= array_access_00037(32 - 16 - 1 downto 0);
  tmp_0019 <= not run_aftrans_Src2In_req_flag_d;
  tmp_0020 <= run_aftrans_Src2In_req_flag and tmp_0019;
  tmp_0021 <= run_aftrans_Src2In_req_flag or run_aftrans_Src2In_req_flag_d;
  tmp_0022 <= run_aftrans_Src2In_req_flag or run_aftrans_Src2In_req_flag_d;
  tmp_0023 <= '1' when binary_expr_00049 = '1' else '0';
  tmp_0024 <= '1' when binary_expr_00049 = '0' else '0';
  tmp_0025 <= '1' when class_m0_0002_fetch_busy = '0' else '0';
  tmp_0026 <= '1' when class_m0_0002_fetch_req = '0' else '0';
  tmp_0027 <= tmp_0025 and tmp_0026;
  tmp_0028 <= '1' when tmp_0027 = '1' else '0';
  tmp_0029 <= '1' when binary_expr_00054 = '1' else '0';
  tmp_0030 <= '1' when binary_expr_00054 = '0' else '0';
  tmp_0031 <= '1' when class_m0_0002_read_busy = '0' else '0';
  tmp_0032 <= '1' when class_m0_0002_read_req = '0' else '0';
  tmp_0033 <= tmp_0031 and tmp_0032;
  tmp_0034 <= '1' when tmp_0033 = '1' else '0';
  tmp_0035 <= '1' when binary_expr_00063 = '1' else '0';
  tmp_0036 <= '1' when binary_expr_00063 = '0' else '0';
  tmp_0037 <= '1' when class_m0_0002_fetch_busy = '0' else '0';
  tmp_0038 <= '1' when class_m0_0002_fetch_req = '0' else '0';
  tmp_0039 <= tmp_0037 and tmp_0038;
  tmp_0040 <= '1' when tmp_0039 = '1' else '0';
  tmp_0041 <= '1' when binary_expr_00068 = '1' else '0';
  tmp_0042 <= '1' when binary_expr_00068 = '0' else '0';
  tmp_0043 <= '1' when class_m0_0002_read_busy = '0' else '0';
  tmp_0044 <= '1' when class_m0_0002_read_req = '0' else '0';
  tmp_0045 <= tmp_0043 and tmp_0044;
  tmp_0046 <= '1' when tmp_0045 = '1' else '0';
  tmp_0047 <= '1' when run_aftrans_Src2In_method /= run_aftrans_Src2In_method_S_0000 else '0';
  tmp_0048 <= '1' when run_aftrans_Src2In_method /= run_aftrans_Src2In_method_S_0001 else '0';
  tmp_0049 <= tmp_0048 and run_aftrans_Src2In_req_flag_edge;
  tmp_0050 <= tmp_0047 and tmp_0049;
  tmp_0051 <= '1' when run_aftrans_Src2In_size_0045 >= class_BS_0006 else '0';
  tmp_0052 <= run_aftrans_Src2In_offset_0048(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0053 <= run_aftrans_Src2In_src_addr_0042 + binary_expr_00051;
  tmp_0054 <= '1' when run_aftrans_Src2In_i_0053 < class_BS_0006 else '0';
  tmp_0055 <= run_aftrans_Src2In_i_0053 + X"00000001";
  tmp_0056 <= run_aftrans_Src2In_offset_0048 + run_aftrans_Src2In_i_0053;
  tmp_0057 <= run_aftrans_Src2In_offset_0048 + class_BS_0006;
  tmp_0058 <= run_aftrans_Src2In_size_0045 - class_BS_0006;
  tmp_0059 <= '1' when run_aftrans_Src2In_size_0045 = X"00000000" else '0';
  tmp_0060 <= run_aftrans_Src2In_offset_0048(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0061 <= run_aftrans_Src2In_src_addr_0042 + binary_expr_00065;
  tmp_0062 <= '1' when run_aftrans_Src2In_i_0067 < run_aftrans_Src2In_size_0045 else '0';
  tmp_0063 <= run_aftrans_Src2In_i_0067 + X"00000001";
  tmp_0064 <= run_aftrans_Src2In_offset_0048 + run_aftrans_Src2In_i_0067;
  tmp_0065 <= not run_aftrans_Src2Cmp_req_flag_d;
  tmp_0066 <= run_aftrans_Src2Cmp_req_flag and tmp_0065;
  tmp_0067 <= run_aftrans_Src2Cmp_req_flag or run_aftrans_Src2Cmp_req_flag_d;
  tmp_0068 <= run_aftrans_Src2Cmp_req_flag or run_aftrans_Src2Cmp_req_flag_d;
  tmp_0069 <= '1' when binary_expr_00082 = '1' else '0';
  tmp_0070 <= '1' when binary_expr_00082 = '0' else '0';
  tmp_0071 <= '1' when binary_expr_00087 = '1' else '0';
  tmp_0072 <= '1' when binary_expr_00087 = '0' else '0';
  tmp_0073 <= '1' when binary_expr_00096 = '1' else '0';
  tmp_0074 <= '1' when binary_expr_00096 = '0' else '0';
  tmp_0075 <= '1' when binary_expr_00101 = '1' else '0';
  tmp_0076 <= '1' when binary_expr_00101 = '0' else '0';
  tmp_0077 <= '1' when run_aftrans_Src2Cmp_method /= run_aftrans_Src2Cmp_method_S_0000 else '0';
  tmp_0078 <= '1' when run_aftrans_Src2Cmp_method /= run_aftrans_Src2Cmp_method_S_0001 else '0';
  tmp_0079 <= tmp_0078 and run_aftrans_Src2Cmp_req_flag_edge;
  tmp_0080 <= tmp_0077 and tmp_0079;
  tmp_0081 <= '1' when run_aftrans_Src2Cmp_size_0078 >= class_BS_0006 else '0';
  tmp_0082 <= run_aftrans_Src2Cmp_offset_0081(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0083 <= run_aftrans_Src2Cmp_src_addr_0075 + binary_expr_00084;
  tmp_0084 <= '1' when run_aftrans_Src2Cmp_i_0086 < class_BS_0006 else '0';
  tmp_0085 <= run_aftrans_Src2Cmp_i_0086 + X"00000001";
  tmp_0086 <= run_aftrans_Src2Cmp_offset_0081 + run_aftrans_Src2Cmp_i_0086;
  tmp_0087 <= run_aftrans_Src2Cmp_offset_0081 + class_BS_0006;
  tmp_0088 <= run_aftrans_Src2Cmp_size_0078 - class_BS_0006;
  tmp_0089 <= '1' when run_aftrans_Src2Cmp_size_0078 = X"00000000" else '0';
  tmp_0090 <= run_aftrans_Src2Cmp_offset_0081(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0091 <= run_aftrans_Src2Cmp_src_addr_0075 + binary_expr_00098;
  tmp_0092 <= '1' when run_aftrans_Src2Cmp_i_0100 < run_aftrans_Src2Cmp_size_0078 else '0';
  tmp_0093 <= run_aftrans_Src2Cmp_i_0100 + X"00000001";
  tmp_0094 <= run_aftrans_Src2Cmp_offset_0081 + run_aftrans_Src2Cmp_i_0100;
  tmp_0095 <= not run_aftrans_Out2Dst_req_flag_d;
  tmp_0096 <= run_aftrans_Out2Dst_req_flag and tmp_0095;
  tmp_0097 <= run_aftrans_Out2Dst_req_flag or run_aftrans_Out2Dst_req_flag_d;
  tmp_0098 <= run_aftrans_Out2Dst_req_flag or run_aftrans_Out2Dst_req_flag_d;
  tmp_0099 <= '1' when binary_expr_00115 = '1' else '0';
  tmp_0100 <= '1' when binary_expr_00115 = '0' else '0';
  tmp_0101 <= '1' when binary_expr_00117 = '1' else '0';
  tmp_0102 <= '1' when binary_expr_00117 = '0' else '0';
  tmp_0103 <= '1' when class_m0_0002_write_busy = '0' else '0';
  tmp_0104 <= '1' when class_m0_0002_write_req = '0' else '0';
  tmp_0105 <= tmp_0103 and tmp_0104;
  tmp_0106 <= '1' when tmp_0105 = '1' else '0';
  tmp_0107 <= '1' when class_m0_0002_flush_busy = '0' else '0';
  tmp_0108 <= '1' when class_m0_0002_flush_req = '0' else '0';
  tmp_0109 <= tmp_0107 and tmp_0108;
  tmp_0110 <= '1' when tmp_0109 = '1' else '0';
  tmp_0111 <= '1' when binary_expr_00129 = '1' else '0';
  tmp_0112 <= '1' when binary_expr_00129 = '0' else '0';
  tmp_0113 <= '1' when binary_expr_00131 = '1' else '0';
  tmp_0114 <= '1' when binary_expr_00131 = '0' else '0';
  tmp_0115 <= '1' when class_m0_0002_write_busy = '0' else '0';
  tmp_0116 <= '1' when class_m0_0002_write_req = '0' else '0';
  tmp_0117 <= tmp_0115 and tmp_0116;
  tmp_0118 <= '1' when tmp_0117 = '1' else '0';
  tmp_0119 <= '1' when class_m0_0002_flush_busy = '0' else '0';
  tmp_0120 <= '1' when class_m0_0002_flush_req = '0' else '0';
  tmp_0121 <= tmp_0119 and tmp_0120;
  tmp_0122 <= '1' when tmp_0121 = '1' else '0';
  tmp_0123 <= '1' when run_aftrans_Out2Dst_method /= run_aftrans_Out2Dst_method_S_0000 else '0';
  tmp_0124 <= '1' when run_aftrans_Out2Dst_method /= run_aftrans_Out2Dst_method_S_0001 else '0';
  tmp_0125 <= tmp_0124 and run_aftrans_Out2Dst_req_flag_edge;
  tmp_0126 <= tmp_0123 and tmp_0125;
  tmp_0127 <= '1' when run_aftrans_Out2Dst_size_0111 >= class_BS_0006 else '0';
  tmp_0128 <= '1' when run_aftrans_Out2Dst_i_0116 < class_BS_0006 else '0';
  tmp_0129 <= run_aftrans_Out2Dst_i_0116 + X"00000001";
  tmp_0130 <= run_aftrans_Out2Dst_offset_0114 + run_aftrans_Out2Dst_i_0116;
  tmp_0131 <= run_aftrans_Out2Dst_offset_0114(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0132 <= run_aftrans_Out2Dst_dst_addr_0108 + binary_expr_00125;
  tmp_0133 <= run_aftrans_Out2Dst_offset_0114 + class_BS_0006;
  tmp_0134 <= run_aftrans_Out2Dst_size_0111 - class_BS_0006;
  tmp_0135 <= '1' when run_aftrans_Out2Dst_size_0111 = X"00000000" else '0';
  tmp_0136 <= '1' when run_aftrans_Out2Dst_i_0130 < run_aftrans_Out2Dst_size_0111 else '0';
  tmp_0137 <= run_aftrans_Out2Dst_i_0130 + X"00000001";
  tmp_0138 <= run_aftrans_Out2Dst_offset_0114 + run_aftrans_Out2Dst_i_0130;
  tmp_0139 <= run_aftrans_Out2Dst_offset_0114(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0140 <= run_aftrans_Out2Dst_dst_addr_0108 + binary_expr_00139;
  tmp_0141 <= not run_memcpy_req_flag_d;
  tmp_0142 <= run_memcpy_req_flag and tmp_0141;
  tmp_0143 <= run_memcpy_req_flag or run_memcpy_req_flag_d;
  tmp_0144 <= run_memcpy_req_flag or run_memcpy_req_flag_d;
  tmp_0145 <= '1' when binary_expr_00151 = '1' else '0';
  tmp_0146 <= '1' when binary_expr_00151 = '0' else '0';
  tmp_0147 <= '1' when class_m0_0002_fetch_busy = '0' else '0';
  tmp_0148 <= '1' when class_m0_0002_fetch_req = '0' else '0';
  tmp_0149 <= tmp_0147 and tmp_0148;
  tmp_0150 <= '1' when tmp_0149 = '1' else '0';
  tmp_0151 <= '1' when class_m0_0002_flush_busy = '0' else '0';
  tmp_0152 <= '1' when class_m0_0002_flush_req = '0' else '0';
  tmp_0153 <= tmp_0151 and tmp_0152;
  tmp_0154 <= '1' when tmp_0153 = '1' else '0';
  tmp_0155 <= '1' when binary_expr_00160 = '1' else '0';
  tmp_0156 <= '1' when binary_expr_00160 = '0' else '0';
  tmp_0157 <= '1' when class_m0_0002_fetch_busy = '0' else '0';
  tmp_0158 <= '1' when class_m0_0002_fetch_req = '0' else '0';
  tmp_0159 <= tmp_0157 and tmp_0158;
  tmp_0160 <= '1' when tmp_0159 = '1' else '0';
  tmp_0161 <= '1' when class_m0_0002_flush_busy = '0' else '0';
  tmp_0162 <= '1' when class_m0_0002_flush_req = '0' else '0';
  tmp_0163 <= tmp_0161 and tmp_0162;
  tmp_0164 <= '1' when tmp_0163 = '1' else '0';
  tmp_0165 <= '1' when run_memcpy_method /= run_memcpy_method_S_0000 else '0';
  tmp_0166 <= '1' when run_memcpy_method /= run_memcpy_method_S_0001 else '0';
  tmp_0167 <= tmp_0166 and run_memcpy_req_flag_edge;
  tmp_0168 <= tmp_0165 and tmp_0167;
  tmp_0169 <= '1' when run_memcpy_size_0147 >= class_BS_0006 else '0';
  tmp_0170 <= run_memcpy_offset_0150(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0171 <= run_memcpy_src_addr_0141 + binary_expr_00153;
  tmp_0172 <= run_memcpy_offset_0150(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0173 <= run_memcpy_dest_addr_0144 + binary_expr_00156;
  tmp_0174 <= run_memcpy_size_0147 - class_BS_0006;
  tmp_0175 <= run_memcpy_offset_0150 + class_BS_0006;
  tmp_0176 <= '1' when run_memcpy_size_0147 = X"00000000" else '0';
  tmp_0177 <= run_memcpy_offset_0150(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0178 <= run_memcpy_src_addr_0141 + binary_expr_00162;
  tmp_0179 <= run_memcpy_offset_0150(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0180 <= run_memcpy_dest_addr_0144 + binary_expr_00165;
  tmp_0181 <= '1' and '1';
  tmp_0182 <= '1' and '0';
  tmp_0183 <= '1' when class_reset_0008 = '1' else '0';
  tmp_0184 <= '1' when class_reset_0008 = '0' else '0';
  tmp_0185 <= class_counter_0007 + X"00000001";
  tmp_0186 <= '1' when binary_expr_00172 = '1' else '0';
  tmp_0187 <= '1' when binary_expr_00172 = '0' else '0';
  tmp_0188 <= '1' when main_cmd_0173 = X"00000010" else '0';
  tmp_0189 <= '1' when main_cmd_0173 = X"00000011" else '0';
  tmp_0190 <= '1' when main_cmd_0173 = X"00000012" else '0';
  tmp_0191 <= '1' when main_cmd_0173 = X"00000018" else '0';
  tmp_0192 <= '1' when main_cmd_0173 = X"00000019" else '0';
  tmp_0193 <= '1' when main_cmd_0173 = X"0000001a" else '0';
  tmp_0194 <= '1' when main_cmd_0173 = X"0000001b" else '0';
  tmp_0195 <= '1' when main_cmd_0173 = X"00000001" else '0';
  tmp_0196 <= '1' when run_memcpy_busy = '0' else '0';
  tmp_0197 <= '1' when run_memcpy_req_local = '0' else '0';
  tmp_0198 <= tmp_0196 and tmp_0197;
  tmp_0199 <= '1' when tmp_0198 = '1' else '0';
  tmp_0200 <= '1' when run_aftrans_proc_busy = '0' else '0';
  tmp_0201 <= '1' when run_aftrans_proc_req_local = '0' else '0';
  tmp_0202 <= tmp_0200 and tmp_0201;
  tmp_0203 <= '1' when tmp_0202 = '1' else '0';
  tmp_0204 <= '1' when run_aftrans_proc_busy = '0' else '0';
  tmp_0205 <= '1' when run_aftrans_proc_req_local = '0' else '0';
  tmp_0206 <= tmp_0204 and tmp_0205;
  tmp_0207 <= '1' when tmp_0206 = '1' else '0';
  tmp_0208 <= '1' when run_aftrans_proc_busy = '0' else '0';
  tmp_0209 <= '1' when run_aftrans_proc_req_local = '0' else '0';
  tmp_0210 <= tmp_0208 and tmp_0209;
  tmp_0211 <= '1' when tmp_0210 = '1' else '0';
  tmp_0212 <= '1' when run_aftrans_proc_busy = '0' else '0';
  tmp_0213 <= '1' when run_aftrans_proc_req_local = '0' else '0';
  tmp_0214 <= tmp_0212 and tmp_0213;
  tmp_0215 <= '1' when tmp_0214 = '1' else '0';
  tmp_0216 <= '1' when run_aftrans_Out2Dst_busy = '0' else '0';
  tmp_0217 <= '1' when run_aftrans_Out2Dst_req_local = '0' else '0';
  tmp_0218 <= tmp_0216 and tmp_0217;
  tmp_0219 <= '1' when tmp_0218 = '1' else '0';
  tmp_0220 <= '1' when run_aftrans_Src2Cmp_busy = '0' else '0';
  tmp_0221 <= '1' when run_aftrans_Src2Cmp_req_local = '0' else '0';
  tmp_0222 <= tmp_0220 and tmp_0221;
  tmp_0223 <= '1' when tmp_0222 = '1' else '0';
  tmp_0224 <= '1' when run_aftrans_Src2In_busy = '0' else '0';
  tmp_0225 <= '1' when run_aftrans_Src2In_req_local = '0' else '0';
  tmp_0226 <= tmp_0224 and tmp_0225;
  tmp_0227 <= '1' when tmp_0226 = '1' else '0';
  tmp_0228 <= '1' when array_access_00171 = X"00000000" else '0';

  -- sequencers
  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_proc_method <= run_aftrans_proc_method_IDLE;
        run_aftrans_proc_method_delay <= (others => '0');
      else
        case (run_aftrans_proc_method) is
          when run_aftrans_proc_method_IDLE => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0000;
          when run_aftrans_proc_method_S_0000 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0001;
          when run_aftrans_proc_method_S_0001 => 
            if tmp_0003 = '1' then
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0002;
            end if;
          when run_aftrans_proc_method_S_0002 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0003;
          when run_aftrans_proc_method_S_0003 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0004;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0004 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0005;
          when run_aftrans_proc_method_S_0005 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0006;
          when run_aftrans_proc_method_S_0006 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0007;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0007 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0008;
          when run_aftrans_proc_method_S_0008 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0009;
          when run_aftrans_proc_method_S_0009 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0010;
          when run_aftrans_proc_method_S_0010 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0011;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0011 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0012;
          when run_aftrans_proc_method_S_0012 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0013;
          when run_aftrans_proc_method_S_0013 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0014;
          when run_aftrans_proc_method_S_0014 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0015;
          when run_aftrans_proc_method_S_0015 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0016;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0016 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0017;
          when run_aftrans_proc_method_S_0017 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0018;
          when run_aftrans_proc_method_S_0018 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0019;
          when run_aftrans_proc_method_S_0019 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0020;
          when run_aftrans_proc_method_S_0020 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0021;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0021 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0022;
          when run_aftrans_proc_method_S_0022 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0023;
          when run_aftrans_proc_method_S_0023 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0024;
          when run_aftrans_proc_method_S_0024 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0025;
          when run_aftrans_proc_method_S_0025 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0026;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0026 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0027;
          when run_aftrans_proc_method_S_0027 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0028;
          when run_aftrans_proc_method_S_0028 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0029;
          when run_aftrans_proc_method_S_0029 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0030;
          when run_aftrans_proc_method_S_0030 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0031;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0031 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0032;
          when run_aftrans_proc_method_S_0032 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0033;
          when run_aftrans_proc_method_S_0033 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0034;
          when run_aftrans_proc_method_S_0034 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0035;
          when run_aftrans_proc_method_S_0035 => 
            if run_aftrans_proc_method_delay >= 2 then
              run_aftrans_proc_method_delay <= (others => '0');
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0036;
            else
              run_aftrans_proc_method_delay <= run_aftrans_proc_method_delay + 1;
            end if;
          when run_aftrans_proc_method_S_0036 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0037;
          when run_aftrans_proc_method_S_0037 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0038;
          when run_aftrans_proc_method_S_0038 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0039;
          when run_aftrans_proc_method_S_0039 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0040;
          when run_aftrans_proc_method_S_0040 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0041;
          when run_aftrans_proc_method_S_0041 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0042;
          when run_aftrans_proc_method_S_0042 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0042_body;
          when run_aftrans_proc_method_S_0043 => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0000;
          when run_aftrans_proc_method_S_0042_body => 
            run_aftrans_proc_method <= run_aftrans_proc_method_S_0042_wait;
          when run_aftrans_proc_method_S_0042_wait => 
            if proc_ext_call_flag_0042 = '1' then
              run_aftrans_proc_method <= run_aftrans_proc_method_S_0043;
            end if;
          when others => null;
        end case;
        run_aftrans_proc_req_flag_d <= run_aftrans_proc_req_flag;
        if (tmp_0009 and tmp_0011) = '1' then
          run_aftrans_proc_method <= run_aftrans_proc_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_method <= run_aftrans_Src2In_method_IDLE;
        run_aftrans_Src2In_method_delay <= (others => '0');
      else
        case (run_aftrans_Src2In_method) is
          when run_aftrans_Src2In_method_IDLE => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0000;
          when run_aftrans_Src2In_method_S_0000 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0001;
          when run_aftrans_Src2In_method_S_0001 => 
            if tmp_0021 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0002;
            end if;
          when run_aftrans_Src2In_method_S_0002 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0003;
          when run_aftrans_Src2In_method_S_0003 => 
            if run_aftrans_Src2In_method_delay >= 2 then
              run_aftrans_Src2In_method_delay <= (others => '0');
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0004;
            else
              run_aftrans_Src2In_method_delay <= run_aftrans_Src2In_method_delay + 1;
            end if;
          when run_aftrans_Src2In_method_S_0004 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0005;
          when run_aftrans_Src2In_method_S_0005 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0006;
          when run_aftrans_Src2In_method_S_0006 => 
            if run_aftrans_Src2In_method_delay >= 2 then
              run_aftrans_Src2In_method_delay <= (others => '0');
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0007;
            else
              run_aftrans_Src2In_method_delay <= run_aftrans_Src2In_method_delay + 1;
            end if;
          when run_aftrans_Src2In_method_S_0007 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0009;
          when run_aftrans_Src2In_method_S_0009 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0010;
          when run_aftrans_Src2In_method_S_0010 => 
            if tmp_0023 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0012;
            elsif tmp_0024 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0011;
            end if;
          when run_aftrans_Src2In_method_S_0011 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0034;
          when run_aftrans_Src2In_method_S_0012 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0013;
          when run_aftrans_Src2In_method_S_0013 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0014;
          when run_aftrans_Src2In_method_S_0014 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0014_body;
          when run_aftrans_Src2In_method_S_0015 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0016;
          when run_aftrans_Src2In_method_S_0016 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0017;
          when run_aftrans_Src2In_method_S_0017 => 
            if tmp_0029 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0022;
            elsif tmp_0030 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0018;
            end if;
          when run_aftrans_Src2In_method_S_0018 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0029;
          when run_aftrans_Src2In_method_S_0019 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0020;
          when run_aftrans_Src2In_method_S_0020 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0021;
          when run_aftrans_Src2In_method_S_0021 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0016;
          when run_aftrans_Src2In_method_S_0022 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0022_body;
          when run_aftrans_Src2In_method_S_0023 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0024;
          when run_aftrans_Src2In_method_S_0024 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0025;
          when run_aftrans_Src2In_method_S_0025 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0026;
          when run_aftrans_Src2In_method_S_0026 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0028;
          when run_aftrans_Src2In_method_S_0028 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0019;
          when run_aftrans_Src2In_method_S_0029 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0030;
          when run_aftrans_Src2In_method_S_0030 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0033;
          when run_aftrans_Src2In_method_S_0033 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0009;
          when run_aftrans_Src2In_method_S_0034 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0035;
          when run_aftrans_Src2In_method_S_0035 => 
            if tmp_0035 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0037;
            elsif tmp_0036 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0036;
            end if;
          when run_aftrans_Src2In_method_S_0036 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0039;
          when run_aftrans_Src2In_method_S_0037 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0000;
          when run_aftrans_Src2In_method_S_0038 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0036;
          when run_aftrans_Src2In_method_S_0039 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0040;
          when run_aftrans_Src2In_method_S_0040 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0041;
          when run_aftrans_Src2In_method_S_0041 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0041_body;
          when run_aftrans_Src2In_method_S_0042 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0043;
          when run_aftrans_Src2In_method_S_0043 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0044;
          when run_aftrans_Src2In_method_S_0044 => 
            if tmp_0041 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0049;
            elsif tmp_0042 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0045;
            end if;
          when run_aftrans_Src2In_method_S_0045 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0056;
          when run_aftrans_Src2In_method_S_0046 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0047;
          when run_aftrans_Src2In_method_S_0047 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0048;
          when run_aftrans_Src2In_method_S_0048 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0043;
          when run_aftrans_Src2In_method_S_0049 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0049_body;
          when run_aftrans_Src2In_method_S_0050 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0051;
          when run_aftrans_Src2In_method_S_0051 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0052;
          when run_aftrans_Src2In_method_S_0052 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0053;
          when run_aftrans_Src2In_method_S_0053 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0055;
          when run_aftrans_Src2In_method_S_0055 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0046;
          when run_aftrans_Src2In_method_S_0056 => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0000;
          when run_aftrans_Src2In_method_S_0014_body => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0014_wait;
          when run_aftrans_Src2In_method_S_0014_wait => 
            if fetch_ext_call_flag_0014 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0015;
            end if;
          when run_aftrans_Src2In_method_S_0022_body => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0022_wait;
          when run_aftrans_Src2In_method_S_0022_wait => 
            if read_ext_call_flag_0022 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0023;
            end if;
          when run_aftrans_Src2In_method_S_0041_body => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0041_wait;
          when run_aftrans_Src2In_method_S_0041_wait => 
            if fetch_ext_call_flag_0041 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0042;
            end if;
          when run_aftrans_Src2In_method_S_0049_body => 
            run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0049_wait;
          when run_aftrans_Src2In_method_S_0049_wait => 
            if read_ext_call_flag_0049 = '1' then
              run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0050;
            end if;
          when others => null;
        end case;
        run_aftrans_Src2In_req_flag_d <= run_aftrans_Src2In_req_flag;
        if (tmp_0047 and tmp_0049) = '1' then
          run_aftrans_Src2In_method <= run_aftrans_Src2In_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_IDLE;
        run_aftrans_Src2Cmp_method_delay <= (others => '0');
      else
        case (run_aftrans_Src2Cmp_method) is
          when run_aftrans_Src2Cmp_method_IDLE => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0000;
          when run_aftrans_Src2Cmp_method_S_0000 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0001;
          when run_aftrans_Src2Cmp_method_S_0001 => 
            if tmp_0067 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0002;
            end if;
          when run_aftrans_Src2Cmp_method_S_0002 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0003;
          when run_aftrans_Src2Cmp_method_S_0003 => 
            if run_aftrans_Src2Cmp_method_delay >= 2 then
              run_aftrans_Src2Cmp_method_delay <= (others => '0');
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0004;
            else
              run_aftrans_Src2Cmp_method_delay <= run_aftrans_Src2Cmp_method_delay + 1;
            end if;
          when run_aftrans_Src2Cmp_method_S_0004 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0005;
          when run_aftrans_Src2Cmp_method_S_0005 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0006;
          when run_aftrans_Src2Cmp_method_S_0006 => 
            if run_aftrans_Src2Cmp_method_delay >= 2 then
              run_aftrans_Src2Cmp_method_delay <= (others => '0');
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0007;
            else
              run_aftrans_Src2Cmp_method_delay <= run_aftrans_Src2Cmp_method_delay + 1;
            end if;
          when run_aftrans_Src2Cmp_method_S_0007 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0009;
          when run_aftrans_Src2Cmp_method_S_0009 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0010;
          when run_aftrans_Src2Cmp_method_S_0010 => 
            if tmp_0069 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0012;
            elsif tmp_0070 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0011;
            end if;
          when run_aftrans_Src2Cmp_method_S_0011 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0034;
          when run_aftrans_Src2Cmp_method_S_0012 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0013;
          when run_aftrans_Src2Cmp_method_S_0013 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0014;
          when run_aftrans_Src2Cmp_method_S_0014 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0014_body;
          when run_aftrans_Src2Cmp_method_S_0015 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0016;
          when run_aftrans_Src2Cmp_method_S_0016 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0017;
          when run_aftrans_Src2Cmp_method_S_0017 => 
            if tmp_0071 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0022;
            elsif tmp_0072 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0018;
            end if;
          when run_aftrans_Src2Cmp_method_S_0018 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0029;
          when run_aftrans_Src2Cmp_method_S_0019 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0020;
          when run_aftrans_Src2Cmp_method_S_0020 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0021;
          when run_aftrans_Src2Cmp_method_S_0021 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0016;
          when run_aftrans_Src2Cmp_method_S_0022 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0022_body;
          when run_aftrans_Src2Cmp_method_S_0023 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0024;
          when run_aftrans_Src2Cmp_method_S_0024 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0025;
          when run_aftrans_Src2Cmp_method_S_0025 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0026;
          when run_aftrans_Src2Cmp_method_S_0026 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0028;
          when run_aftrans_Src2Cmp_method_S_0028 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0019;
          when run_aftrans_Src2Cmp_method_S_0029 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0030;
          when run_aftrans_Src2Cmp_method_S_0030 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0033;
          when run_aftrans_Src2Cmp_method_S_0033 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0009;
          when run_aftrans_Src2Cmp_method_S_0034 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0035;
          when run_aftrans_Src2Cmp_method_S_0035 => 
            if tmp_0073 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0037;
            elsif tmp_0074 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0036;
            end if;
          when run_aftrans_Src2Cmp_method_S_0036 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0039;
          when run_aftrans_Src2Cmp_method_S_0037 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0000;
          when run_aftrans_Src2Cmp_method_S_0038 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0036;
          when run_aftrans_Src2Cmp_method_S_0039 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0040;
          when run_aftrans_Src2Cmp_method_S_0040 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0041;
          when run_aftrans_Src2Cmp_method_S_0041 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0041_body;
          when run_aftrans_Src2Cmp_method_S_0042 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0043;
          when run_aftrans_Src2Cmp_method_S_0043 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0044;
          when run_aftrans_Src2Cmp_method_S_0044 => 
            if tmp_0075 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0049;
            elsif tmp_0076 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0045;
            end if;
          when run_aftrans_Src2Cmp_method_S_0045 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0056;
          when run_aftrans_Src2Cmp_method_S_0046 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0047;
          when run_aftrans_Src2Cmp_method_S_0047 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0048;
          when run_aftrans_Src2Cmp_method_S_0048 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0043;
          when run_aftrans_Src2Cmp_method_S_0049 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0049_body;
          when run_aftrans_Src2Cmp_method_S_0050 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0051;
          when run_aftrans_Src2Cmp_method_S_0051 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0052;
          when run_aftrans_Src2Cmp_method_S_0052 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0053;
          when run_aftrans_Src2Cmp_method_S_0053 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0055;
          when run_aftrans_Src2Cmp_method_S_0055 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0046;
          when run_aftrans_Src2Cmp_method_S_0056 => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0000;
          when run_aftrans_Src2Cmp_method_S_0014_body => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0014_wait;
          when run_aftrans_Src2Cmp_method_S_0014_wait => 
            if fetch_ext_call_flag_0014 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0015;
            end if;
          when run_aftrans_Src2Cmp_method_S_0022_body => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0022_wait;
          when run_aftrans_Src2Cmp_method_S_0022_wait => 
            if read_ext_call_flag_0022 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0023;
            end if;
          when run_aftrans_Src2Cmp_method_S_0041_body => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0041_wait;
          when run_aftrans_Src2Cmp_method_S_0041_wait => 
            if fetch_ext_call_flag_0041 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0042;
            end if;
          when run_aftrans_Src2Cmp_method_S_0049_body => 
            run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0049_wait;
          when run_aftrans_Src2Cmp_method_S_0049_wait => 
            if read_ext_call_flag_0049 = '1' then
              run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0050;
            end if;
          when others => null;
        end case;
        run_aftrans_Src2Cmp_req_flag_d <= run_aftrans_Src2Cmp_req_flag;
        if (tmp_0077 and tmp_0079) = '1' then
          run_aftrans_Src2Cmp_method <= run_aftrans_Src2Cmp_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_IDLE;
        run_aftrans_Out2Dst_method_delay <= (others => '0');
      else
        case (run_aftrans_Out2Dst_method) is
          when run_aftrans_Out2Dst_method_IDLE => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0000;
          when run_aftrans_Out2Dst_method_S_0000 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0001;
          when run_aftrans_Out2Dst_method_S_0001 => 
            if tmp_0097 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0002;
            end if;
          when run_aftrans_Out2Dst_method_S_0002 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0003;
          when run_aftrans_Out2Dst_method_S_0003 => 
            if run_aftrans_Out2Dst_method_delay >= 2 then
              run_aftrans_Out2Dst_method_delay <= (others => '0');
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0004;
            else
              run_aftrans_Out2Dst_method_delay <= run_aftrans_Out2Dst_method_delay + 1;
            end if;
          when run_aftrans_Out2Dst_method_S_0004 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0005;
          when run_aftrans_Out2Dst_method_S_0005 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0006;
          when run_aftrans_Out2Dst_method_S_0006 => 
            if run_aftrans_Out2Dst_method_delay >= 2 then
              run_aftrans_Out2Dst_method_delay <= (others => '0');
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0007;
            else
              run_aftrans_Out2Dst_method_delay <= run_aftrans_Out2Dst_method_delay + 1;
            end if;
          when run_aftrans_Out2Dst_method_S_0007 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0009;
          when run_aftrans_Out2Dst_method_S_0009 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0010;
          when run_aftrans_Out2Dst_method_S_0010 => 
            if tmp_0099 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0012;
            elsif tmp_0100 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0011;
            end if;
          when run_aftrans_Out2Dst_method_S_0011 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0033;
          when run_aftrans_Out2Dst_method_S_0012 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0013;
          when run_aftrans_Out2Dst_method_S_0013 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0014;
          when run_aftrans_Out2Dst_method_S_0014 => 
            if tmp_0101 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0019;
            elsif tmp_0102 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0015;
            end if;
          when run_aftrans_Out2Dst_method_S_0015 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0025;
          when run_aftrans_Out2Dst_method_S_0016 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0017;
          when run_aftrans_Out2Dst_method_S_0017 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0018;
          when run_aftrans_Out2Dst_method_S_0018 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0013;
          when run_aftrans_Out2Dst_method_S_0019 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0020;
          when run_aftrans_Out2Dst_method_S_0020 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0021;
          when run_aftrans_Out2Dst_method_S_0021 => 
            if run_aftrans_Out2Dst_method_delay >= 2 then
              run_aftrans_Out2Dst_method_delay <= (others => '0');
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0022;
            else
              run_aftrans_Out2Dst_method_delay <= run_aftrans_Out2Dst_method_delay + 1;
            end if;
          when run_aftrans_Out2Dst_method_S_0022 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0023;
          when run_aftrans_Out2Dst_method_S_0023 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0023_body;
          when run_aftrans_Out2Dst_method_S_0024 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0016;
          when run_aftrans_Out2Dst_method_S_0025 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0026;
          when run_aftrans_Out2Dst_method_S_0026 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0027;
          when run_aftrans_Out2Dst_method_S_0027 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0027_body;
          when run_aftrans_Out2Dst_method_S_0028 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0029;
          when run_aftrans_Out2Dst_method_S_0029 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0032;
          when run_aftrans_Out2Dst_method_S_0032 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0009;
          when run_aftrans_Out2Dst_method_S_0033 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0034;
          when run_aftrans_Out2Dst_method_S_0034 => 
            if tmp_0111 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0036;
            elsif tmp_0112 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0035;
            end if;
          when run_aftrans_Out2Dst_method_S_0035 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0038;
          when run_aftrans_Out2Dst_method_S_0036 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0000;
          when run_aftrans_Out2Dst_method_S_0037 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0035;
          when run_aftrans_Out2Dst_method_S_0038 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0039;
          when run_aftrans_Out2Dst_method_S_0039 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0040;
          when run_aftrans_Out2Dst_method_S_0040 => 
            if tmp_0113 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0045;
            elsif tmp_0114 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0041;
            end if;
          when run_aftrans_Out2Dst_method_S_0041 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0051;
          when run_aftrans_Out2Dst_method_S_0042 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0043;
          when run_aftrans_Out2Dst_method_S_0043 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0044;
          when run_aftrans_Out2Dst_method_S_0044 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0039;
          when run_aftrans_Out2Dst_method_S_0045 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0046;
          when run_aftrans_Out2Dst_method_S_0046 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0047;
          when run_aftrans_Out2Dst_method_S_0047 => 
            if run_aftrans_Out2Dst_method_delay >= 2 then
              run_aftrans_Out2Dst_method_delay <= (others => '0');
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0048;
            else
              run_aftrans_Out2Dst_method_delay <= run_aftrans_Out2Dst_method_delay + 1;
            end if;
          when run_aftrans_Out2Dst_method_S_0048 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0049;
          when run_aftrans_Out2Dst_method_S_0049 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0049_body;
          when run_aftrans_Out2Dst_method_S_0050 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0042;
          when run_aftrans_Out2Dst_method_S_0051 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0052;
          when run_aftrans_Out2Dst_method_S_0052 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0053;
          when run_aftrans_Out2Dst_method_S_0053 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0053_body;
          when run_aftrans_Out2Dst_method_S_0054 => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0000;
          when run_aftrans_Out2Dst_method_S_0023_body => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0023_wait;
          when run_aftrans_Out2Dst_method_S_0023_wait => 
            if write_ext_call_flag_0023 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0024;
            end if;
          when run_aftrans_Out2Dst_method_S_0027_body => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0027_wait;
          when run_aftrans_Out2Dst_method_S_0027_wait => 
            if flush_ext_call_flag_0027 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0028;
            end if;
          when run_aftrans_Out2Dst_method_S_0049_body => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0049_wait;
          when run_aftrans_Out2Dst_method_S_0049_wait => 
            if write_ext_call_flag_0049 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0050;
            end if;
          when run_aftrans_Out2Dst_method_S_0053_body => 
            run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0053_wait;
          when run_aftrans_Out2Dst_method_S_0053_wait => 
            if flush_ext_call_flag_0053 = '1' then
              run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0054;
            end if;
          when others => null;
        end case;
        run_aftrans_Out2Dst_req_flag_d <= run_aftrans_Out2Dst_req_flag;
        if (tmp_0123 and tmp_0125) = '1' then
          run_aftrans_Out2Dst_method <= run_aftrans_Out2Dst_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_memcpy_method <= run_memcpy_method_IDLE;
        run_memcpy_method_delay <= (others => '0');
      else
        case (run_memcpy_method) is
          when run_memcpy_method_IDLE => 
            run_memcpy_method <= run_memcpy_method_S_0000;
          when run_memcpy_method_S_0000 => 
            run_memcpy_method <= run_memcpy_method_S_0001;
          when run_memcpy_method_S_0001 => 
            if tmp_0143 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0002;
            end if;
          when run_memcpy_method_S_0002 => 
            run_memcpy_method <= run_memcpy_method_S_0003;
          when run_memcpy_method_S_0003 => 
            if run_memcpy_method_delay >= 2 then
              run_memcpy_method_delay <= (others => '0');
              run_memcpy_method <= run_memcpy_method_S_0004;
            else
              run_memcpy_method_delay <= run_memcpy_method_delay + 1;
            end if;
          when run_memcpy_method_S_0004 => 
            run_memcpy_method <= run_memcpy_method_S_0005;
          when run_memcpy_method_S_0005 => 
            run_memcpy_method <= run_memcpy_method_S_0006;
          when run_memcpy_method_S_0006 => 
            if run_memcpy_method_delay >= 2 then
              run_memcpy_method_delay <= (others => '0');
              run_memcpy_method <= run_memcpy_method_S_0007;
            else
              run_memcpy_method_delay <= run_memcpy_method_delay + 1;
            end if;
          when run_memcpy_method_S_0007 => 
            run_memcpy_method <= run_memcpy_method_S_0008;
          when run_memcpy_method_S_0008 => 
            run_memcpy_method <= run_memcpy_method_S_0009;
          when run_memcpy_method_S_0009 => 
            if run_memcpy_method_delay >= 2 then
              run_memcpy_method_delay <= (others => '0');
              run_memcpy_method <= run_memcpy_method_S_0010;
            else
              run_memcpy_method_delay <= run_memcpy_method_delay + 1;
            end if;
          when run_memcpy_method_S_0010 => 
            run_memcpy_method <= run_memcpy_method_S_0012;
          when run_memcpy_method_S_0012 => 
            run_memcpy_method <= run_memcpy_method_S_0013;
          when run_memcpy_method_S_0013 => 
            if tmp_0145 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0015;
            elsif tmp_0146 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0014;
            end if;
          when run_memcpy_method_S_0014 => 
            run_memcpy_method <= run_memcpy_method_S_0026;
          when run_memcpy_method_S_0015 => 
            run_memcpy_method <= run_memcpy_method_S_0016;
          when run_memcpy_method_S_0016 => 
            run_memcpy_method <= run_memcpy_method_S_0017;
          when run_memcpy_method_S_0017 => 
            run_memcpy_method <= run_memcpy_method_S_0017_body;
          when run_memcpy_method_S_0018 => 
            run_memcpy_method <= run_memcpy_method_S_0019;
          when run_memcpy_method_S_0019 => 
            run_memcpy_method <= run_memcpy_method_S_0020;
          when run_memcpy_method_S_0020 => 
            run_memcpy_method <= run_memcpy_method_S_0020_body;
          when run_memcpy_method_S_0021 => 
            run_memcpy_method <= run_memcpy_method_S_0022;
          when run_memcpy_method_S_0022 => 
            run_memcpy_method <= run_memcpy_method_S_0025;
          when run_memcpy_method_S_0025 => 
            run_memcpy_method <= run_memcpy_method_S_0012;
          when run_memcpy_method_S_0026 => 
            run_memcpy_method <= run_memcpy_method_S_0027;
          when run_memcpy_method_S_0027 => 
            if tmp_0155 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0029;
            elsif tmp_0156 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0028;
            end if;
          when run_memcpy_method_S_0028 => 
            run_memcpy_method <= run_memcpy_method_S_0031;
          when run_memcpy_method_S_0029 => 
            run_memcpy_method <= run_memcpy_method_S_0000;
          when run_memcpy_method_S_0030 => 
            run_memcpy_method <= run_memcpy_method_S_0028;
          when run_memcpy_method_S_0031 => 
            run_memcpy_method <= run_memcpy_method_S_0032;
          when run_memcpy_method_S_0032 => 
            run_memcpy_method <= run_memcpy_method_S_0033;
          when run_memcpy_method_S_0033 => 
            run_memcpy_method <= run_memcpy_method_S_0033_body;
          when run_memcpy_method_S_0034 => 
            run_memcpy_method <= run_memcpy_method_S_0035;
          when run_memcpy_method_S_0035 => 
            run_memcpy_method <= run_memcpy_method_S_0036;
          when run_memcpy_method_S_0036 => 
            run_memcpy_method <= run_memcpy_method_S_0036_body;
          when run_memcpy_method_S_0037 => 
            run_memcpy_method <= run_memcpy_method_S_0000;
          when run_memcpy_method_S_0017_body => 
            run_memcpy_method <= run_memcpy_method_S_0017_wait;
          when run_memcpy_method_S_0017_wait => 
            if fetch_ext_call_flag_0017 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0018;
            end if;
          when run_memcpy_method_S_0020_body => 
            run_memcpy_method <= run_memcpy_method_S_0020_wait;
          when run_memcpy_method_S_0020_wait => 
            if flush_ext_call_flag_0020 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0021;
            end if;
          when run_memcpy_method_S_0033_body => 
            run_memcpy_method <= run_memcpy_method_S_0033_wait;
          when run_memcpy_method_S_0033_wait => 
            if fetch_ext_call_flag_0033 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0034;
            end if;
          when run_memcpy_method_S_0036_body => 
            run_memcpy_method <= run_memcpy_method_S_0036_wait;
          when run_memcpy_method_S_0036_wait => 
            if flush_ext_call_flag_0036 = '1' then
              run_memcpy_method <= run_memcpy_method_S_0037;
            end if;
          when others => null;
        end case;
        run_memcpy_req_flag_d <= run_memcpy_req_flag;
        if (tmp_0165 and tmp_0167) = '1' then
          run_memcpy_method <= run_memcpy_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        clock_method <= clock_method_IDLE;
        clock_method_delay <= (others => '0');
      else
        case (clock_method) is
          when clock_method_IDLE => 
            clock_method <= clock_method_S_0000;
          when clock_method_S_0000 => 
            clock_method <= clock_method_S_0001;
          when clock_method_S_0001 => 
            clock_method <= clock_method_S_0002;
          when clock_method_S_0002 => 
            if tmp_0181 = '1' then
              clock_method <= clock_method_S_0004;
            elsif tmp_0182 = '1' then
              clock_method <= clock_method_S_0003;
            end if;
          when clock_method_S_0003 => 
            clock_method <= clock_method_S_0013;
          when clock_method_S_0004 => 
            if tmp_0183 = '1' then
              clock_method <= clock_method_S_0006;
            elsif tmp_0184 = '1' then
              clock_method <= clock_method_S_0009;
            end if;
          when clock_method_S_0005 => 
            clock_method <= clock_method_S_0012;
          when clock_method_S_0006 => 
            clock_method <= clock_method_S_0008;
          when clock_method_S_0008 => 
            clock_method <= clock_method_S_0005;
          when clock_method_S_0009 => 
            clock_method <= clock_method_S_0010;
          when clock_method_S_0010 => 
            clock_method <= clock_method_S_0011;
          when clock_method_S_0011 => 
            clock_method <= clock_method_S_0005;
          when clock_method_S_0012 => 
            clock_method <= clock_method_S_0002;
          when clock_method_S_0013 => 
            clock_method <= clock_method_S_0000;
          when others => null;
        end case;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        main_method <= main_method_IDLE;
        main_method_delay <= (others => '0');
      else
        case (main_method) is
          when main_method_IDLE => 
            main_method <= main_method_S_0000;
          when main_method_S_0000 => 
            main_method <= main_method_S_0001;
          when main_method_S_0001 => 
            main_method <= main_method_S_0002;
          when main_method_S_0002 => 
            main_method <= main_method_S_0003;
          when main_method_S_0003 => 
            main_method <= main_method_S_0005;
          when main_method_S_0005 => 
            main_method <= main_method_S_0006;
          when main_method_S_0006 => 
            if main_method_delay >= 2 then
              main_method_delay <= (others => '0');
              main_method <= main_method_S_0007;
            else
              main_method_delay <= main_method_delay + 1;
            end if;
          when main_method_S_0007 => 
            main_method <= main_method_S_0008;
          when main_method_S_0008 => 
            if tmp_0186 = '1' then
              main_method <= main_method_S_0010;
            elsif tmp_0187 = '1' then
              main_method <= main_method_S_0009;
            end if;
          when main_method_S_0009 => 
            main_method <= main_method_S_0011;
          when main_method_S_0010 => 
            main_method <= main_method_S_0005;
          when main_method_S_0011 => 
            main_method <= main_method_S_0012;
          when main_method_S_0012 => 
            if main_method_delay >= 2 then
              main_method_delay <= (others => '0');
              main_method <= main_method_S_0013;
            else
              main_method_delay <= main_method_delay + 1;
            end if;
          when main_method_S_0013 => 
            main_method <= main_method_S_0015;
          when main_method_S_0015 => 
            if tmp_0188 = '1' then
              main_method <= main_method_S_0063;
            elsif tmp_0189 = '1' then
              main_method <= main_method_S_0060;
            elsif tmp_0190 = '1' then
              main_method <= main_method_S_0057;
            elsif tmp_0191 = '1' then
              main_method <= main_method_S_0046;
            elsif tmp_0192 = '1' then
              main_method <= main_method_S_0035;
            elsif tmp_0193 = '1' then
              main_method <= main_method_S_0028;
            elsif tmp_0194 = '1' then
              main_method <= main_method_S_0021;
            elsif tmp_0195 = '1' then
              main_method <= main_method_S_0018;
            else
              main_method <= main_method_S_0017;
            end if;
          when main_method_S_0016 => 
            main_method <= main_method_S_0066;
          when main_method_S_0017 => 
            main_method <= main_method_S_0016;
          when main_method_S_0018 => 
            main_method <= main_method_S_0018_body;
          when main_method_S_0019 => 
            main_method <= main_method_S_0016;
          when main_method_S_0020 => 
            main_method <= main_method_S_0017;
          when main_method_S_0021 => 
            main_method <= main_method_S_0022;
          when main_method_S_0022 => 
            main_method <= main_method_S_0023;
          when main_method_S_0023 => 
            main_method <= main_method_S_0024;
          when main_method_S_0024 => 
            main_method <= main_method_S_0025;
          when main_method_S_0025 => 
            main_method <= main_method_S_0025_body;
          when main_method_S_0026 => 
            main_method <= main_method_S_0016;
          when main_method_S_0027 => 
            main_method <= main_method_S_0018;
          when main_method_S_0028 => 
            main_method <= main_method_S_0029;
          when main_method_S_0029 => 
            main_method <= main_method_S_0030;
          when main_method_S_0030 => 
            main_method <= main_method_S_0031;
          when main_method_S_0031 => 
            main_method <= main_method_S_0032;
          when main_method_S_0032 => 
            main_method <= main_method_S_0032_body;
          when main_method_S_0033 => 
            main_method <= main_method_S_0016;
          when main_method_S_0034 => 
            main_method <= main_method_S_0021;
          when main_method_S_0035 => 
            main_method <= main_method_S_0036;
          when main_method_S_0036 => 
            main_method <= main_method_S_0037;
          when main_method_S_0037 => 
            main_method <= main_method_S_0038;
          when main_method_S_0038 => 
            main_method <= main_method_S_0039;
          when main_method_S_0039 => 
            main_method <= main_method_S_0039_body;
          when main_method_S_0040 => 
            main_method <= main_method_S_0041;
          when main_method_S_0041 => 
            main_method <= main_method_S_0042;
          when main_method_S_0042 => 
            main_method <= main_method_S_0043;
          when main_method_S_0043 => 
            main_method <= main_method_S_0044;
          when main_method_S_0044 => 
            main_method <= main_method_S_0016;
          when main_method_S_0045 => 
            main_method <= main_method_S_0028;
          when main_method_S_0046 => 
            main_method <= main_method_S_0047;
          when main_method_S_0047 => 
            main_method <= main_method_S_0048;
          when main_method_S_0048 => 
            main_method <= main_method_S_0049;
          when main_method_S_0049 => 
            main_method <= main_method_S_0050;
          when main_method_S_0050 => 
            main_method <= main_method_S_0050_body;
          when main_method_S_0051 => 
            main_method <= main_method_S_0052;
          when main_method_S_0052 => 
            main_method <= main_method_S_0053;
          when main_method_S_0053 => 
            main_method <= main_method_S_0054;
          when main_method_S_0054 => 
            main_method <= main_method_S_0055;
          when main_method_S_0055 => 
            main_method <= main_method_S_0016;
          when main_method_S_0056 => 
            main_method <= main_method_S_0035;
          when main_method_S_0057 => 
            main_method <= main_method_S_0057_body;
          when main_method_S_0058 => 
            main_method <= main_method_S_0016;
          when main_method_S_0059 => 
            main_method <= main_method_S_0046;
          when main_method_S_0060 => 
            main_method <= main_method_S_0060_body;
          when main_method_S_0061 => 
            main_method <= main_method_S_0016;
          when main_method_S_0062 => 
            main_method <= main_method_S_0057;
          when main_method_S_0063 => 
            main_method <= main_method_S_0063_body;
          when main_method_S_0064 => 
            main_method <= main_method_S_0016;
          when main_method_S_0065 => 
            main_method <= main_method_S_0060;
          when main_method_S_0066 => 
            main_method <= main_method_S_0067;
          when main_method_S_0067 => 
            main_method <= main_method_S_0069;
          when main_method_S_0069 => 
            main_method <= main_method_S_0070;
          when main_method_S_0070 => 
            main_method <= main_method_S_0072;
          when main_method_S_0072 => 
            main_method <= main_method_S_0000;
          when main_method_S_0018_body => 
            main_method <= main_method_S_0018_wait;
          when main_method_S_0018_wait => 
            if run_memcpy_call_flag_0018 = '1' then
              main_method <= main_method_S_0019;
            end if;
          when main_method_S_0025_body => 
            main_method <= main_method_S_0025_wait;
          when main_method_S_0025_wait => 
            if run_aftrans_proc_call_flag_0025 = '1' then
              main_method <= main_method_S_0026;
            end if;
          when main_method_S_0032_body => 
            main_method <= main_method_S_0032_wait;
          when main_method_S_0032_wait => 
            if run_aftrans_proc_call_flag_0032 = '1' then
              main_method <= main_method_S_0033;
            end if;
          when main_method_S_0039_body => 
            main_method <= main_method_S_0039_wait;
          when main_method_S_0039_wait => 
            if run_aftrans_proc_call_flag_0039 = '1' then
              main_method <= main_method_S_0040;
            end if;
          when main_method_S_0050_body => 
            main_method <= main_method_S_0050_wait;
          when main_method_S_0050_wait => 
            if run_aftrans_proc_call_flag_0050 = '1' then
              main_method <= main_method_S_0051;
            end if;
          when main_method_S_0057_body => 
            main_method <= main_method_S_0057_wait;
          when main_method_S_0057_wait => 
            if run_aftrans_Out2Dst_call_flag_0057 = '1' then
              main_method <= main_method_S_0058;
            end if;
          when main_method_S_0060_body => 
            main_method <= main_method_S_0060_wait;
          when main_method_S_0060_wait => 
            if run_aftrans_Src2Cmp_call_flag_0060 = '1' then
              main_method <= main_method_S_0061;
            end if;
          when main_method_S_0063_body => 
            main_method <= main_method_S_0063_wait;
          when main_method_S_0063_wait => 
            if run_aftrans_Src2In_call_flag_0063 = '1' then
              main_method <= main_method_S_0064;
            end if;
          when others => null;
        end case;
      end if;
    end if;
  end process;


  class_s0_0000_clk <= clk_sig;

  class_s0_0000_reset <= reset_sig;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_s0_0000_data_address <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0003 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000001";
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0006 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000002";
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0010 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000003";
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0015 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000004";
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0020 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000005";
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0025 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000006";
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0030 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000007";
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0035 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_address <= X"00000008";
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0003 and run_aftrans_Src2In_method_delay = 0 then
          class_s0_0000_data_address <= X"00000001";
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0006 and run_aftrans_Src2In_method_delay = 0 then
          class_s0_0000_data_address <= X"00000002";
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0003 and run_aftrans_Src2Cmp_method_delay = 0 then
          class_s0_0000_data_address <= X"00000001";
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0006 and run_aftrans_Src2Cmp_method_delay = 0 then
          class_s0_0000_data_address <= X"00000002";
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0003 and run_aftrans_Out2Dst_method_delay = 0 then
          class_s0_0000_data_address <= X"00000001";
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0006 and run_aftrans_Out2Dst_method_delay = 0 then
          class_s0_0000_data_address <= X"00000002";
        elsif run_memcpy_method = run_memcpy_method_S_0003 and run_memcpy_method_delay = 0 then
          class_s0_0000_data_address <= X"00000001";
        elsif run_memcpy_method = run_memcpy_method_S_0006 and run_memcpy_method_delay = 0 then
          class_s0_0000_data_address <= X"00000002";
        elsif run_memcpy_method = run_memcpy_method_S_0009 and run_memcpy_method_delay = 0 then
          class_s0_0000_data_address <= X"00000003";
        elsif main_method = main_method_S_0003 then
          class_s0_0000_data_address <= X"00000000";
        elsif main_method = main_method_S_0006 and main_method_delay = 0 then
          class_s0_0000_data_address <= X"00000000";
        elsif main_method = main_method_S_0012 and main_method_delay = 0 then
          class_s0_0000_data_address <= X"00000000";
        elsif main_method = main_method_S_0041 then
          class_s0_0000_data_address <= X"00000002";
        elsif main_method = main_method_S_0052 then
          class_s0_0000_data_address <= X"00000002";
        elsif main_method = main_method_S_0067 then
          class_s0_0000_data_address <= X"00000001";
        elsif main_method = main_method_S_0070 then
          class_s0_0000_data_address <= X"00000000";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_s0_0000_data_din <= (others => '0');
      else
        if main_method = main_method_S_0003 then
          class_s0_0000_data_din <= X"00000000";
        elsif main_method = main_method_S_0043 then
          class_s0_0000_data_din <= std_logic_vector(field_access_00188);
        elsif main_method = main_method_S_0054 then
          class_s0_0000_data_din <= std_logic_vector(field_access_00194);
        elsif main_method = main_method_S_0067 then
          class_s0_0000_data_din <= std_logic_vector(class_counter_0007);
        elsif main_method = main_method_S_0070 then
          class_s0_0000_data_din <= X"00000000";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_s0_0000_data_we <= '0';
      else
        if main_method = main_method_S_0003 then
          class_s0_0000_data_we <= '1';
        elsif main_method = main_method_S_0043 then
          class_s0_0000_data_we <= '1';
        elsif main_method = main_method_S_0054 then
          class_s0_0000_data_we <= '1';
        elsif main_method = main_method_S_0067 then
          class_s0_0000_data_we <= '1';
        elsif main_method = main_method_S_0070 then
          class_s0_0000_data_we <= '1';
        else
          class_s0_0000_data_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_s0_0000_data_oe <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0003 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0006 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0010 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0015 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0020 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0025 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0030 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0035 and run_aftrans_proc_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0003 and run_aftrans_Src2In_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0006 and run_aftrans_Src2In_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0003 and run_aftrans_Src2Cmp_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0006 and run_aftrans_Src2Cmp_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0003 and run_aftrans_Out2Dst_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0006 and run_aftrans_Out2Dst_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_memcpy_method = run_memcpy_method_S_0003 and run_memcpy_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_memcpy_method = run_memcpy_method_S_0006 and run_memcpy_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif run_memcpy_method = run_memcpy_method_S_0009 and run_memcpy_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif main_method = main_method_S_0006 and main_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        elsif main_method = main_method_S_0012 and main_method_delay = 0 then
          class_s0_0000_data_oe <= '1';
        else
          class_s0_0000_data_oe <= '0';
        end if;
      end if;
    end if;
  end process;

  class_s0_0000_axi_reader_ARADDR <= class_s0_0000_axi_reader_ARADDR_exp_sig;

  class_s0_0000_axi_reader_ARVALID <= class_s0_0000_axi_reader_ARVALID_exp_sig;

  class_s0_0000_axi_reader_RREADY <= class_s0_0000_axi_reader_RREADY_exp_sig;

  class_s0_0000_axi_writer_AWADDR <= class_s0_0000_axi_writer_AWADDR_exp_sig;

  class_s0_0000_axi_writer_AWVALID <= class_s0_0000_axi_writer_AWVALID_exp_sig;

  class_s0_0000_axi_writer_WDATA <= class_s0_0000_axi_writer_WDATA_exp_sig;

  class_s0_0000_axi_writer_WVALID <= class_s0_0000_axi_writer_WVALID_exp_sig;

  class_s0_0000_axi_writer_WSTRB <= class_s0_0000_axi_writer_WSTRB_exp_sig;

  class_s0_0000_axi_writer_BREADY <= class_s0_0000_axi_writer_BREADY_exp_sig;

  class_m0_0002_clk <= clk_sig;

  class_m0_0002_reset <= reset_sig;

  class_m0_0002_class_obj_0000_forbid_exp <= class_m0_0002_class_obj_0000_forbid_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp <= class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_reader_RDATA_exp <= class_m0_0002_class_obj_0000_axi_reader_RDATA_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_reader_RRESP_exp <= class_m0_0002_class_obj_0000_axi_reader_RRESP_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_reader_RLAST_exp <= class_m0_0002_class_obj_0000_axi_reader_RLAST_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_reader_RVALID_exp <= class_m0_0002_class_obj_0000_axi_reader_RVALID_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp <= class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_writer_WREADY_exp <= class_m0_0002_class_obj_0000_axi_writer_WREADY_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_writer_BRESP_exp <= class_m0_0002_class_obj_0000_axi_writer_BRESP_exp_exp_sig;

  class_m0_0002_class_obj_0000_axi_writer_BVALID_exp <= class_m0_0002_class_obj_0000_axi_writer_BVALID_exp_exp_sig;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_flush_addr <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0027_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_flush_addr <= binary_expr_00126;
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0053_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_flush_addr <= binary_expr_00140;
        elsif run_memcpy_method = run_memcpy_method_S_0020_body and run_memcpy_method_delay = 0 then
          class_m0_0002_flush_addr <= binary_expr_00157;
        elsif run_memcpy_method = run_memcpy_method_S_0036_body and run_memcpy_method_delay = 0 then
          class_m0_0002_flush_addr <= binary_expr_00166;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_flush_burst <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0027_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_flush_burst <= class_BS_0006;
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0053_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_flush_burst <= run_aftrans_Out2Dst_size_0111;
        elsif run_memcpy_method = run_memcpy_method_S_0020_body and run_memcpy_method_delay = 0 then
          class_m0_0002_flush_burst <= class_BS_0006;
        elsif run_memcpy_method = run_memcpy_method_S_0036_body and run_memcpy_method_delay = 0 then
          class_m0_0002_flush_burst <= run_memcpy_size_0147;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_fetch_addr <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0014_body and run_aftrans_Src2In_method_delay = 0 then
          class_m0_0002_fetch_addr <= binary_expr_00052;
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0041_body and run_aftrans_Src2In_method_delay = 0 then
          class_m0_0002_fetch_addr <= binary_expr_00066;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0014_body and run_aftrans_Src2Cmp_method_delay = 0 then
          class_m0_0002_fetch_addr <= binary_expr_00085;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0041_body and run_aftrans_Src2Cmp_method_delay = 0 then
          class_m0_0002_fetch_addr <= binary_expr_00099;
        elsif run_memcpy_method = run_memcpy_method_S_0017_body and run_memcpy_method_delay = 0 then
          class_m0_0002_fetch_addr <= binary_expr_00154;
        elsif run_memcpy_method = run_memcpy_method_S_0033_body and run_memcpy_method_delay = 0 then
          class_m0_0002_fetch_addr <= binary_expr_00163;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_fetch_burst <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0014_body and run_aftrans_Src2In_method_delay = 0 then
          class_m0_0002_fetch_burst <= class_BS_0006;
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0041_body and run_aftrans_Src2In_method_delay = 0 then
          class_m0_0002_fetch_burst <= run_aftrans_Src2In_size_0045;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0014_body and run_aftrans_Src2Cmp_method_delay = 0 then
          class_m0_0002_fetch_burst <= class_BS_0006;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0041_body and run_aftrans_Src2Cmp_method_delay = 0 then
          class_m0_0002_fetch_burst <= run_aftrans_Src2Cmp_size_0078;
        elsif run_memcpy_method = run_memcpy_method_S_0017_body and run_memcpy_method_delay = 0 then
          class_m0_0002_fetch_burst <= class_BS_0006;
        elsif run_memcpy_method = run_memcpy_method_S_0033_body and run_memcpy_method_delay = 0 then
          class_m0_0002_fetch_burst <= run_memcpy_size_0147;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_read_offset <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0022_body and run_aftrans_Src2In_method_delay = 0 then
          class_m0_0002_read_offset <= run_aftrans_Src2In_i_0053;
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0049_body and run_aftrans_Src2In_method_delay = 0 then
          class_m0_0002_read_offset <= run_aftrans_Src2In_i_0067;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0022_body and run_aftrans_Src2Cmp_method_delay = 0 then
          class_m0_0002_read_offset <= run_aftrans_Src2Cmp_i_0086;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0049_body and run_aftrans_Src2Cmp_method_delay = 0 then
          class_m0_0002_read_offset <= run_aftrans_Src2Cmp_i_0100;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_write_offset <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0023_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_write_offset <= run_aftrans_Out2Dst_i_0116;
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0049_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_write_offset <= run_aftrans_Out2Dst_i_0130;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_write_data <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0023_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_write_data <= run_aftrans_Out2Dst_d_0119;
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0049_body and run_aftrans_Out2Dst_method_delay = 0 then
          class_m0_0002_write_data <= run_aftrans_Out2Dst_d_0133;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_flush_req <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0027_body then
          class_m0_0002_flush_req <= '1';
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0053_body then
          class_m0_0002_flush_req <= '1';
        elsif run_memcpy_method = run_memcpy_method_S_0020_body then
          class_m0_0002_flush_req <= '1';
        elsif run_memcpy_method = run_memcpy_method_S_0036_body then
          class_m0_0002_flush_req <= '1';
        else
          class_m0_0002_flush_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_fetch_req <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0014_body then
          class_m0_0002_fetch_req <= '1';
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0041_body then
          class_m0_0002_fetch_req <= '1';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0014_body then
          class_m0_0002_fetch_req <= '1';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0041_body then
          class_m0_0002_fetch_req <= '1';
        elsif run_memcpy_method = run_memcpy_method_S_0017_body then
          class_m0_0002_fetch_req <= '1';
        elsif run_memcpy_method = run_memcpy_method_S_0033_body then
          class_m0_0002_fetch_req <= '1';
        else
          class_m0_0002_fetch_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_read_req <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0022_body then
          class_m0_0002_read_req <= '1';
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0049_body then
          class_m0_0002_read_req <= '1';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0022_body then
          class_m0_0002_read_req <= '1';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0049_body then
          class_m0_0002_read_req <= '1';
        else
          class_m0_0002_read_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_m0_0002_write_req <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0023_body then
          class_m0_0002_write_req <= '1';
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0049_body then
          class_m0_0002_write_req <= '1';
        else
          class_m0_0002_write_req <= '0';
        end if;
      end if;
    end if;
  end process;

  class_at_0004_clk <= clk_sig;

  class_at_0004_reset <= reset_sig;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_width_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0039 then
          class_at_0004_width_in <= run_aftrans_proc_width_0009;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_width_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0039 then
          class_at_0004_width_we <= '1';
        else
          class_at_0004_width_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_height_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0041 then
          class_at_0004_height_in <= run_aftrans_proc_height_0012;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_height_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0041 then
          class_at_0004_height_we <= '1';
        else
          class_at_0004_height_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_inData_address <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0026 then
          class_at_0004_inData_address <= binary_expr_00059;
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0053 then
          class_at_0004_inData_address <= binary_expr_00073;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_inData_we <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0026 then
          class_at_0004_inData_we <= '1';
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0053 then
          class_at_0004_inData_we <= '1';
        else
          class_at_0004_inData_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_inData_din <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0026 then
          class_at_0004_inData_din <= run_aftrans_Src2In_d_0056;
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0053 then
          class_at_0004_inData_din <= run_aftrans_Src2In_d_0070;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_outData_address <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0021 and run_aftrans_Out2Dst_method_delay = 0 then
          class_at_0004_outData_address <= binary_expr_00121;
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0047 and run_aftrans_Out2Dst_method_delay = 0 then
          class_at_0004_outData_address <= binary_expr_00135;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_outData_oe <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0021 and run_aftrans_Out2Dst_method_delay = 0 then
          class_at_0004_outData_oe <= '1';
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0047 and run_aftrans_Out2Dst_method_delay = 0 then
          class_at_0004_outData_oe <= '1';
        else
          class_at_0004_outData_oe <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_cmpData_address <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0026 then
          class_at_0004_cmpData_address <= binary_expr_00092;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0053 then
          class_at_0004_cmpData_address <= binary_expr_00106;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_cmpData_we <= '0';
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0026 then
          class_at_0004_cmpData_we <= '1';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0053 then
          class_at_0004_cmpData_we <= '1';
        else
          class_at_0004_cmpData_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_cmpData_din <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0026 then
          class_at_0004_cmpData_din <= run_aftrans_Src2Cmp_d_0089;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0053 then
          class_at_0004_cmpData_din <= run_aftrans_Src2Cmp_d_0103;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat00_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0012 then
          class_at_0004_mat00_in <= cast_expr_00018;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat00_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0012 then
          class_at_0004_mat00_we <= '1';
        else
          class_at_0004_mat00_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat01_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0017 then
          class_at_0004_mat01_in <= cast_expr_00022;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat01_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0017 then
          class_at_0004_mat01_we <= '1';
        else
          class_at_0004_mat01_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat02_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0022 then
          class_at_0004_mat02_in <= cast_expr_00026;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat02_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0022 then
          class_at_0004_mat02_we <= '1';
        else
          class_at_0004_mat02_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat10_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0027 then
          class_at_0004_mat10_in <= cast_expr_00030;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat10_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0027 then
          class_at_0004_mat10_we <= '1';
        else
          class_at_0004_mat10_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat11_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0032 then
          class_at_0004_mat11_in <= cast_expr_00034;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat11_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0032 then
          class_at_0004_mat11_we <= '1';
        else
          class_at_0004_mat11_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat12_in <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0037 then
          class_at_0004_mat12_in <= cast_expr_00038;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_mat12_we <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0037 then
          class_at_0004_mat12_we <= '1';
        else
          class_at_0004_mat12_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_modeInterpolation_in <= '0';
      else
        if main_method = main_method_S_0022 then
          class_at_0004_modeInterpolation_in <= '0';
        elsif main_method = main_method_S_0029 then
          class_at_0004_modeInterpolation_in <= '1';
        elsif main_method = main_method_S_0036 then
          class_at_0004_modeInterpolation_in <= '0';
        elsif main_method = main_method_S_0047 then
          class_at_0004_modeInterpolation_in <= '1';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_modeInterpolation_we <= '0';
      else
        if main_method = main_method_S_0022 then
          class_at_0004_modeInterpolation_we <= '1';
        elsif main_method = main_method_S_0029 then
          class_at_0004_modeInterpolation_we <= '1';
        elsif main_method = main_method_S_0036 then
          class_at_0004_modeInterpolation_we <= '1';
        elsif main_method = main_method_S_0047 then
          class_at_0004_modeInterpolation_we <= '1';
        else
          class_at_0004_modeInterpolation_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_modeCompare_in <= '0';
      else
        if main_method = main_method_S_0024 then
          class_at_0004_modeCompare_in <= '0';
        elsif main_method = main_method_S_0031 then
          class_at_0004_modeCompare_in <= '0';
        elsif main_method = main_method_S_0038 then
          class_at_0004_modeCompare_in <= '1';
        elsif main_method = main_method_S_0049 then
          class_at_0004_modeCompare_in <= '1';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_modeCompare_we <= '0';
      else
        if main_method = main_method_S_0024 then
          class_at_0004_modeCompare_we <= '1';
        elsif main_method = main_method_S_0031 then
          class_at_0004_modeCompare_we <= '1';
        elsif main_method = main_method_S_0038 then
          class_at_0004_modeCompare_we <= '1';
        elsif main_method = main_method_S_0049 then
          class_at_0004_modeCompare_we <= '1';
        else
          class_at_0004_modeCompare_we <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_at_0004_proc_req <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0042_body then
          class_at_0004_proc_req <= '1';
        else
          class_at_0004_proc_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_counter_0007 <= X"00000000";
      else
        if clock_method = clock_method_S_0006 then
          class_counter_0007 <= X"00000000";
        elsif clock_method = clock_method_S_0010 then
          class_counter_0007 <= unary_expr_00167;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_reset_0008 <= '1';
      else
        if clock_method = clock_method_S_0006 then
          class_reset_0008 <= '0';
        elsif main_method = main_method_S_0013 then
          class_reset_0008 <= '1';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_proc_width_0009 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0004 then
          run_aftrans_proc_width_0009 <= array_access_00011;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00011 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0003 and run_aftrans_proc_method_delay = 2 then
          array_access_00011 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_proc_height_0012 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0007 then
          run_aftrans_proc_height_0012 <= array_access_00014;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00014 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0006 and run_aftrans_proc_method_delay = 2 then
          array_access_00014 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00015 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0008 then
          field_access_00015 <= class_at_0004_mat00_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00017 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0010 and run_aftrans_proc_method_delay = 2 then
          array_access_00017 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00018 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0011 then
          cast_expr_00018 <= tmp_0013;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00019 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0013 then
          field_access_00019 <= class_at_0004_mat01_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00021 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0015 and run_aftrans_proc_method_delay = 2 then
          array_access_00021 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00022 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0016 then
          cast_expr_00022 <= tmp_0014;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00023 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0018 then
          field_access_00023 <= class_at_0004_mat02_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00025 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0020 and run_aftrans_proc_method_delay = 2 then
          array_access_00025 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00026 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0021 then
          cast_expr_00026 <= tmp_0015;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00027 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0023 then
          field_access_00027 <= class_at_0004_mat10_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00029 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0025 and run_aftrans_proc_method_delay = 2 then
          array_access_00029 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00030 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0026 then
          cast_expr_00030 <= tmp_0016;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00031 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0028 then
          field_access_00031 <= class_at_0004_mat11_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00033 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0030 and run_aftrans_proc_method_delay = 2 then
          array_access_00033 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00034 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0031 then
          cast_expr_00034 <= tmp_0017;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00035 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0033 then
          field_access_00035 <= class_at_0004_mat12_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00037 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0035 and run_aftrans_proc_method_delay = 2 then
          array_access_00037 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00038 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0036 then
          cast_expr_00038 <= tmp_0018;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00039 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0038 then
          field_access_00039 <= class_at_0004_width_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00040 <= (others => '0');
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0040 then
          field_access_00040 <= class_at_0004_height_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_src_addr_0042 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0004 then
          run_aftrans_Src2In_src_addr_0042 <= array_access_00044;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00044 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0003 and run_aftrans_Src2In_method_delay = 2 then
          array_access_00044 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_size_0045 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0007 then
          run_aftrans_Src2In_size_0045 <= array_access_00047;
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0030 then
          run_aftrans_Src2In_size_0045 <= binary_expr_00062;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00047 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0006 and run_aftrans_Src2In_method_delay = 2 then
          array_access_00047 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_offset_0048 <= X"00000000";
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0007 then
          run_aftrans_Src2In_offset_0048 <= X"00000000";
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0030 then
          run_aftrans_Src2In_offset_0048 <= binary_expr_00061;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00049 <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0009 then
          binary_expr_00049 <= tmp_0051;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00063 <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0034 then
          binary_expr_00063 <= tmp_0059;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00065 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0039 then
          binary_expr_00065 <= tmp_0060;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00066 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0040 then
          binary_expr_00066 <= tmp_0061;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00051 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0012 then
          binary_expr_00051 <= tmp_0052;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00052 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0013 then
          binary_expr_00052 <= tmp_0053;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00061 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0029 then
          binary_expr_00061 <= tmp_0057;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00062 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0029 then
          binary_expr_00062 <= tmp_0058;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_i_0053 <= X"00000000";
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0015 then
          run_aftrans_Src2In_i_0053 <= X"00000000";
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0020 then
          run_aftrans_Src2In_i_0053 <= unary_expr_00055;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00054 <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0016 then
          binary_expr_00054 <= tmp_0054;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00055 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0019 then
          unary_expr_00055 <= tmp_0055;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_d_0056 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0023 then
          run_aftrans_Src2In_d_0056 <= method_result_00057;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00057 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0022_wait then
          method_result_00057 <= class_m0_0002_read_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00059 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0025 then
          binary_expr_00059 <= tmp_0056;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_i_0067 <= X"00000000";
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0042 then
          run_aftrans_Src2In_i_0067 <= X"00000000";
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0047 then
          run_aftrans_Src2In_i_0067 <= unary_expr_00069;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00068 <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0043 then
          binary_expr_00068 <= tmp_0062;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00069 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0046 then
          unary_expr_00069 <= tmp_0063;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_d_0070 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0050 then
          run_aftrans_Src2In_d_0070 <= method_result_00071;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00071 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0049_wait then
          method_result_00071 <= class_m0_0002_read_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00073 <= (others => '0');
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0052 then
          binary_expr_00073 <= tmp_0064;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_src_addr_0075 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0004 then
          run_aftrans_Src2Cmp_src_addr_0075 <= array_access_00077;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00077 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0003 and run_aftrans_Src2Cmp_method_delay = 2 then
          array_access_00077 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_size_0078 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0007 then
          run_aftrans_Src2Cmp_size_0078 <= array_access_00080;
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0030 then
          run_aftrans_Src2Cmp_size_0078 <= binary_expr_00095;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00080 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0006 and run_aftrans_Src2Cmp_method_delay = 2 then
          array_access_00080 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_offset_0081 <= X"00000000";
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0007 then
          run_aftrans_Src2Cmp_offset_0081 <= X"00000000";
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0030 then
          run_aftrans_Src2Cmp_offset_0081 <= binary_expr_00094;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00082 <= '0';
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0009 then
          binary_expr_00082 <= tmp_0081;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00096 <= '0';
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0034 then
          binary_expr_00096 <= tmp_0089;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00098 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0039 then
          binary_expr_00098 <= tmp_0090;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00099 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0040 then
          binary_expr_00099 <= tmp_0091;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00084 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0012 then
          binary_expr_00084 <= tmp_0082;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00085 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0013 then
          binary_expr_00085 <= tmp_0083;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00094 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0029 then
          binary_expr_00094 <= tmp_0087;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00095 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0029 then
          binary_expr_00095 <= tmp_0088;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_i_0086 <= X"00000000";
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0015 then
          run_aftrans_Src2Cmp_i_0086 <= X"00000000";
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0020 then
          run_aftrans_Src2Cmp_i_0086 <= unary_expr_00088;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00087 <= '0';
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0016 then
          binary_expr_00087 <= tmp_0084;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00088 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0019 then
          unary_expr_00088 <= tmp_0085;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_d_0089 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0023 then
          run_aftrans_Src2Cmp_d_0089 <= method_result_00090;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00090 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0022_wait then
          method_result_00090 <= class_m0_0002_read_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00092 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0025 then
          binary_expr_00092 <= tmp_0086;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_i_0100 <= X"00000000";
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0042 then
          run_aftrans_Src2Cmp_i_0100 <= X"00000000";
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0047 then
          run_aftrans_Src2Cmp_i_0100 <= unary_expr_00102;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00101 <= '0';
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0043 then
          binary_expr_00101 <= tmp_0092;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00102 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0046 then
          unary_expr_00102 <= tmp_0093;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_d_0103 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0050 then
          run_aftrans_Src2Cmp_d_0103 <= method_result_00104;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00104 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0049_wait then
          method_result_00104 <= class_m0_0002_read_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00106 <= (others => '0');
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0052 then
          binary_expr_00106 <= tmp_0094;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_dst_addr_0108 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0004 then
          run_aftrans_Out2Dst_dst_addr_0108 <= array_access_00110;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00110 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0003 and run_aftrans_Out2Dst_method_delay = 2 then
          array_access_00110 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_size_0111 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0007 then
          run_aftrans_Out2Dst_size_0111 <= array_access_00113;
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0029 then
          run_aftrans_Out2Dst_size_0111 <= binary_expr_00128;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00113 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0006 and run_aftrans_Out2Dst_method_delay = 2 then
          array_access_00113 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_offset_0114 <= X"00000000";
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0007 then
          run_aftrans_Out2Dst_offset_0114 <= X"00000000";
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0029 then
          run_aftrans_Out2Dst_offset_0114 <= binary_expr_00127;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00115 <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0009 then
          binary_expr_00115 <= tmp_0127;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00129 <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0033 then
          binary_expr_00129 <= tmp_0135;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00139 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0051 then
          binary_expr_00139 <= tmp_0139;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00140 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0052 then
          binary_expr_00140 <= tmp_0140;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00125 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0025 then
          binary_expr_00125 <= tmp_0131;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00126 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0026 then
          binary_expr_00126 <= tmp_0132;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00127 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0028 then
          binary_expr_00127 <= tmp_0133;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00128 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0028 then
          binary_expr_00128 <= tmp_0134;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_i_0116 <= X"00000000";
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0012 then
          run_aftrans_Out2Dst_i_0116 <= X"00000000";
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0017 then
          run_aftrans_Out2Dst_i_0116 <= unary_expr_00118;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00117 <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0013 then
          binary_expr_00117 <= tmp_0128;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00118 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0016 then
          unary_expr_00118 <= tmp_0129;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_d_0119 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0022 then
          run_aftrans_Out2Dst_d_0119 <= array_access_00122;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00121 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0020 then
          binary_expr_00121 <= tmp_0130;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00122 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0021 and run_aftrans_Out2Dst_method_delay = 2 then
          array_access_00122 <= class_at_0004_outData_dout;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_i_0130 <= X"00000000";
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0038 then
          run_aftrans_Out2Dst_i_0130 <= X"00000000";
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0043 then
          run_aftrans_Out2Dst_i_0130 <= unary_expr_00132;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00131 <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0039 then
          binary_expr_00131 <= tmp_0136;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00132 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0042 then
          unary_expr_00132 <= tmp_0137;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_d_0133 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0048 then
          run_aftrans_Out2Dst_d_0133 <= array_access_00136;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00135 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0046 then
          binary_expr_00135 <= tmp_0138;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00136 <= (others => '0');
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0047 and run_aftrans_Out2Dst_method_delay = 2 then
          array_access_00136 <= class_at_0004_outData_dout;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_memcpy_src_addr_0141 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0004 then
          run_memcpy_src_addr_0141 <= array_access_00143;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00143 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0003 and run_memcpy_method_delay = 2 then
          array_access_00143 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_memcpy_dest_addr_0144 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0007 then
          run_memcpy_dest_addr_0144 <= array_access_00146;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00146 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0006 and run_memcpy_method_delay = 2 then
          array_access_00146 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_memcpy_size_0147 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0010 then
          run_memcpy_size_0147 <= array_access_00149;
        elsif run_memcpy_method = run_memcpy_method_S_0022 then
          run_memcpy_size_0147 <= binary_expr_00158;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00149 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0009 and run_memcpy_method_delay = 2 then
          array_access_00149 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_memcpy_offset_0150 <= X"00000000";
      else
        if run_memcpy_method = run_memcpy_method_S_0010 then
          run_memcpy_offset_0150 <= X"00000000";
        elsif run_memcpy_method = run_memcpy_method_S_0022 then
          run_memcpy_offset_0150 <= binary_expr_00159;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00151 <= '0';
      else
        if run_memcpy_method = run_memcpy_method_S_0012 then
          binary_expr_00151 <= tmp_0169;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00160 <= '0';
      else
        if run_memcpy_method = run_memcpy_method_S_0026 then
          binary_expr_00160 <= tmp_0176;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00162 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0031 then
          binary_expr_00162 <= tmp_0177;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00163 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0032 then
          binary_expr_00163 <= tmp_0178;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00165 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0034 then
          binary_expr_00165 <= tmp_0179;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00166 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0035 then
          binary_expr_00166 <= tmp_0180;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00153 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0015 then
          binary_expr_00153 <= tmp_0170;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00154 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0016 then
          binary_expr_00154 <= tmp_0171;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00156 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0018 then
          binary_expr_00156 <= tmp_0172;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00157 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0019 then
          binary_expr_00157 <= tmp_0173;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00158 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0021 then
          binary_expr_00158 <= tmp_0174;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00159 <= (others => '0');
      else
        if run_memcpy_method = run_memcpy_method_S_0021 then
          binary_expr_00159 <= tmp_0175;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00167 <= (others => '0');
      else
        if clock_method = clock_method_S_0009 then
          unary_expr_00167 <= tmp_0185;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00171 <= (others => '0');
      else
        if main_method = main_method_S_0006 and main_method_delay = 2 then
          array_access_00171 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00172 <= '0';
      else
        if main_method = main_method_S_0007 then
          binary_expr_00172 <= tmp_0228;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        main_cmd_0173 <= (others => '0');
      else
        if main_method = main_method_S_0013 then
          main_cmd_0173 <= array_access_00175;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00175 <= (others => '0');
      else
        if main_method = main_method_S_0012 and main_method_delay = 2 then
          array_access_00175 <= signed(class_s0_0000_data_dout);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00177 <= '0';
      else
        if main_method = main_method_S_0021 then
          field_access_00177 <= class_at_0004_modeInterpolation_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00178 <= '0';
      else
        if main_method = main_method_S_0023 then
          field_access_00178 <= class_at_0004_modeCompare_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00180 <= '0';
      else
        if main_method = main_method_S_0028 then
          field_access_00180 <= class_at_0004_modeInterpolation_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00181 <= '0';
      else
        if main_method = main_method_S_0030 then
          field_access_00181 <= class_at_0004_modeCompare_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00183 <= '0';
      else
        if main_method = main_method_S_0035 then
          field_access_00183 <= class_at_0004_modeInterpolation_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00184 <= '0';
      else
        if main_method = main_method_S_0037 then
          field_access_00184 <= class_at_0004_modeCompare_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00188 <= (others => '0');
      else
        if main_method = main_method_S_0042 then
          field_access_00188 <= class_at_0004_diffCompare_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00189 <= '0';
      else
        if main_method = main_method_S_0046 then
          field_access_00189 <= class_at_0004_modeInterpolation_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00190 <= '0';
      else
        if main_method = main_method_S_0048 then
          field_access_00190 <= class_at_0004_modeCompare_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00194 <= (others => '0');
      else
        if main_method = main_method_S_0053 then
          field_access_00194 <= class_at_0004_diffCompare_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_proc_busy <= '0';
      else
        if run_aftrans_proc_method = run_aftrans_proc_method_S_0000 then
          run_aftrans_proc_busy <= '0';
        elsif run_aftrans_proc_method = run_aftrans_proc_method_S_0001 then
          run_aftrans_proc_busy <= tmp_0004;
        end if;
      end if;
    end if;
  end process;

  run_aftrans_proc_req_flag <= run_aftrans_proc_req_local;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_proc_req_local <= '0';
      else
        if main_method = main_method_S_0025_body then
          run_aftrans_proc_req_local <= '1';
        elsif main_method = main_method_S_0032_body then
          run_aftrans_proc_req_local <= '1';
        elsif main_method = main_method_S_0039_body then
          run_aftrans_proc_req_local <= '1';
        elsif main_method = main_method_S_0050_body then
          run_aftrans_proc_req_local <= '1';
        else
          run_aftrans_proc_req_local <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_busy <= '0';
      else
        if run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0000 then
          run_aftrans_Src2In_busy <= '0';
        elsif run_aftrans_Src2In_method = run_aftrans_Src2In_method_S_0001 then
          run_aftrans_Src2In_busy <= tmp_0022;
        end if;
      end if;
    end if;
  end process;

  run_aftrans_Src2In_req_flag <= run_aftrans_Src2In_req_local;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2In_req_local <= '0';
      else
        if main_method = main_method_S_0063_body then
          run_aftrans_Src2In_req_local <= '1';
        else
          run_aftrans_Src2In_req_local <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_busy <= '0';
      else
        if run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0000 then
          run_aftrans_Src2Cmp_busy <= '0';
        elsif run_aftrans_Src2Cmp_method = run_aftrans_Src2Cmp_method_S_0001 then
          run_aftrans_Src2Cmp_busy <= tmp_0068;
        end if;
      end if;
    end if;
  end process;

  run_aftrans_Src2Cmp_req_flag <= run_aftrans_Src2Cmp_req_local;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Src2Cmp_req_local <= '0';
      else
        if main_method = main_method_S_0060_body then
          run_aftrans_Src2Cmp_req_local <= '1';
        else
          run_aftrans_Src2Cmp_req_local <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_busy <= '0';
      else
        if run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0000 then
          run_aftrans_Out2Dst_busy <= '0';
        elsif run_aftrans_Out2Dst_method = run_aftrans_Out2Dst_method_S_0001 then
          run_aftrans_Out2Dst_busy <= tmp_0098;
        end if;
      end if;
    end if;
  end process;

  run_aftrans_Out2Dst_req_flag <= run_aftrans_Out2Dst_req_local;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_aftrans_Out2Dst_req_local <= '0';
      else
        if main_method = main_method_S_0057_body then
          run_aftrans_Out2Dst_req_local <= '1';
        else
          run_aftrans_Out2Dst_req_local <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_memcpy_busy <= '0';
      else
        if run_memcpy_method = run_memcpy_method_S_0000 then
          run_memcpy_busy <= '0';
        elsif run_memcpy_method = run_memcpy_method_S_0001 then
          run_memcpy_busy <= tmp_0144;
        end if;
      end if;
    end if;
  end process;

  run_memcpy_req_flag <= run_memcpy_req_local;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        run_memcpy_req_local <= '0';
      else
        if main_method = main_method_S_0018_body then
          run_memcpy_req_local <= '1';
        else
          run_memcpy_req_local <= '0';
        end if;
      end if;
    end if;
  end process;

  run_aftrans_proc_req_flag_edge <= tmp_0002;

  proc_ext_call_flag_0042 <= tmp_0008;

  run_aftrans_Src2In_req_flag_edge <= tmp_0020;

  fetch_ext_call_flag_0014 <= tmp_0028;

  read_ext_call_flag_0022 <= tmp_0034;

  fetch_ext_call_flag_0041 <= tmp_0040;

  read_ext_call_flag_0049 <= tmp_0046;

  run_aftrans_Src2Cmp_req_flag_edge <= tmp_0066;

  run_aftrans_Out2Dst_req_flag_edge <= tmp_0096;

  write_ext_call_flag_0023 <= tmp_0106;

  flush_ext_call_flag_0027 <= tmp_0110;

  write_ext_call_flag_0049 <= tmp_0118;

  flush_ext_call_flag_0053 <= tmp_0122;

  run_memcpy_req_flag_edge <= tmp_0142;

  fetch_ext_call_flag_0017 <= tmp_0150;

  flush_ext_call_flag_0020 <= tmp_0154;

  fetch_ext_call_flag_0033 <= tmp_0160;

  flush_ext_call_flag_0036 <= tmp_0164;

  run_memcpy_call_flag_0018 <= tmp_0199;

  run_aftrans_proc_call_flag_0025 <= tmp_0203;

  run_aftrans_proc_call_flag_0032 <= tmp_0207;

  run_aftrans_proc_call_flag_0039 <= tmp_0211;

  run_aftrans_proc_call_flag_0050 <= tmp_0215;

  run_aftrans_Out2Dst_call_flag_0057 <= tmp_0219;

  run_aftrans_Src2Cmp_call_flag_0060 <= tmp_0223;

  run_aftrans_Src2In_call_flag_0063 <= tmp_0227;


  inst_class_s0_0000 : axi_lite_slave_32
  port map(
    clk => class_s0_0000_clk,
    reset => class_s0_0000_reset,
    data_length => class_s0_0000_data_length,
    data_address => class_s0_0000_data_address,
    data_din => class_s0_0000_data_din,
    data_dout => class_s0_0000_data_dout,
    data_we => class_s0_0000_data_we,
    data_oe => class_s0_0000_data_oe,
    axi_reader_ARADDR => class_s0_0000_axi_reader_ARADDR,
    axi_reader_ARVALID => class_s0_0000_axi_reader_ARVALID,
    axi_reader_ARREADY => class_s0_0000_axi_reader_ARREADY,
    axi_reader_RDATA => class_s0_0000_axi_reader_RDATA,
    axi_reader_RRESP => class_s0_0000_axi_reader_RRESP,
    axi_reader_RVALID => class_s0_0000_axi_reader_RVALID,
    axi_reader_RREADY => class_s0_0000_axi_reader_RREADY,
    axi_writer_AWADDR => class_s0_0000_axi_writer_AWADDR,
    axi_writer_AWVALID => class_s0_0000_axi_writer_AWVALID,
    axi_writer_AWREADY => class_s0_0000_axi_writer_AWREADY,
    axi_writer_WDATA => class_s0_0000_axi_writer_WDATA,
    axi_writer_WVALID => class_s0_0000_axi_writer_WVALID,
    axi_writer_WREADY => class_s0_0000_axi_writer_WREADY,
    axi_writer_WSTRB => class_s0_0000_axi_writer_WSTRB,
    axi_writer_BRESP => class_s0_0000_axi_writer_BRESP,
    axi_writer_BVALID => class_s0_0000_axi_writer_BVALID,
    axi_writer_BREADY => class_s0_0000_axi_writer_BREADY
  );

  inst_class_m0_0002 : synthesijer_lib_axi_AXIMemIface32RTLTest
  port map(
    clk => class_m0_0002_clk,
    reset => class_m0_0002_reset,
    class_obj_0000_forbid_exp => class_m0_0002_class_obj_0000_forbid_exp,
    class_obj_0000_axi_reader_ARADDR_exp => class_m0_0002_class_obj_0000_axi_reader_ARADDR_exp,
    class_obj_0000_axi_reader_ARLEN_exp => class_m0_0002_class_obj_0000_axi_reader_ARLEN_exp,
    class_obj_0000_axi_reader_ARVALID_exp => class_m0_0002_class_obj_0000_axi_reader_ARVALID_exp,
    class_obj_0000_axi_reader_ARREADY_exp => class_m0_0002_class_obj_0000_axi_reader_ARREADY_exp,
    class_obj_0000_axi_reader_ARSIZE_exp => class_m0_0002_class_obj_0000_axi_reader_ARSIZE_exp,
    class_obj_0000_axi_reader_ARBURST_exp => class_m0_0002_class_obj_0000_axi_reader_ARBURST_exp,
    class_obj_0000_axi_reader_ARCACHE_exp => class_m0_0002_class_obj_0000_axi_reader_ARCACHE_exp,
    class_obj_0000_axi_reader_ARPROT_exp => class_m0_0002_class_obj_0000_axi_reader_ARPROT_exp,
    class_obj_0000_axi_reader_RDATA_exp => class_m0_0002_class_obj_0000_axi_reader_RDATA_exp,
    class_obj_0000_axi_reader_RRESP_exp => class_m0_0002_class_obj_0000_axi_reader_RRESP_exp,
    class_obj_0000_axi_reader_RLAST_exp => class_m0_0002_class_obj_0000_axi_reader_RLAST_exp,
    class_obj_0000_axi_reader_RVALID_exp => class_m0_0002_class_obj_0000_axi_reader_RVALID_exp,
    class_obj_0000_axi_reader_RREADY_exp => class_m0_0002_class_obj_0000_axi_reader_RREADY_exp,
    class_obj_0000_axi_writer_AWADDR_exp => class_m0_0002_class_obj_0000_axi_writer_AWADDR_exp,
    class_obj_0000_axi_writer_AWLEN_exp => class_m0_0002_class_obj_0000_axi_writer_AWLEN_exp,
    class_obj_0000_axi_writer_AWVALID_exp => class_m0_0002_class_obj_0000_axi_writer_AWVALID_exp,
    class_obj_0000_axi_writer_AWSIZE_exp => class_m0_0002_class_obj_0000_axi_writer_AWSIZE_exp,
    class_obj_0000_axi_writer_AWBURST_exp => class_m0_0002_class_obj_0000_axi_writer_AWBURST_exp,
    class_obj_0000_axi_writer_AWCACHE_exp => class_m0_0002_class_obj_0000_axi_writer_AWCACHE_exp,
    class_obj_0000_axi_writer_AWPROT_exp => class_m0_0002_class_obj_0000_axi_writer_AWPROT_exp,
    class_obj_0000_axi_writer_AWREADY_exp => class_m0_0002_class_obj_0000_axi_writer_AWREADY_exp,
    class_obj_0000_axi_writer_WDATA_exp => class_m0_0002_class_obj_0000_axi_writer_WDATA_exp,
    class_obj_0000_axi_writer_WLAST_exp => class_m0_0002_class_obj_0000_axi_writer_WLAST_exp,
    class_obj_0000_axi_writer_WVALID_exp => class_m0_0002_class_obj_0000_axi_writer_WVALID_exp,
    class_obj_0000_axi_writer_WREADY_exp => class_m0_0002_class_obj_0000_axi_writer_WREADY_exp,
    class_obj_0000_axi_writer_WSTRB_exp => class_m0_0002_class_obj_0000_axi_writer_WSTRB_exp,
    class_obj_0000_axi_writer_BRESP_exp => class_m0_0002_class_obj_0000_axi_writer_BRESP_exp,
    class_obj_0000_axi_writer_BVALID_exp => class_m0_0002_class_obj_0000_axi_writer_BVALID_exp,
    class_obj_0000_axi_writer_BREADY_exp => class_m0_0002_class_obj_0000_axi_writer_BREADY_exp,
    flush_addr => class_m0_0002_flush_addr,
    flush_burst => class_m0_0002_flush_burst,
    fetch_addr => class_m0_0002_fetch_addr,
    fetch_burst => class_m0_0002_fetch_burst,
    read_offset => class_m0_0002_read_offset,
    write_offset => class_m0_0002_write_offset,
    write_data => class_m0_0002_write_data,
    flush_busy => class_m0_0002_flush_busy,
    flush_req => class_m0_0002_flush_req,
    fetch_busy => class_m0_0002_fetch_busy,
    fetch_req => class_m0_0002_fetch_req,
    read_return => class_m0_0002_read_return,
    read_busy => class_m0_0002_read_busy,
    read_req => class_m0_0002_read_req,
    write_busy => class_m0_0002_write_busy,
    write_req => class_m0_0002_write_req
  );

  inst_class_at_0004 : AffineTransform
  port map(
    clk => class_at_0004_clk,
    reset => class_at_0004_reset,
    width_in => class_at_0004_width_in,
    width_we => class_at_0004_width_we,
    width_out => class_at_0004_width_out,
    height_in => class_at_0004_height_in,
    height_we => class_at_0004_height_we,
    height_out => class_at_0004_height_out,
    inData_address => class_at_0004_inData_address,
    inData_we => class_at_0004_inData_we,
    inData_oe => class_at_0004_inData_oe,
    inData_din => class_at_0004_inData_din,
    inData_dout => class_at_0004_inData_dout,
    inData_length => class_at_0004_inData_length,
    outData_address => class_at_0004_outData_address,
    outData_we => class_at_0004_outData_we,
    outData_oe => class_at_0004_outData_oe,
    outData_din => class_at_0004_outData_din,
    outData_dout => class_at_0004_outData_dout,
    outData_length => class_at_0004_outData_length,
    cmpData_address => class_at_0004_cmpData_address,
    cmpData_we => class_at_0004_cmpData_we,
    cmpData_oe => class_at_0004_cmpData_oe,
    cmpData_din => class_at_0004_cmpData_din,
    cmpData_dout => class_at_0004_cmpData_dout,
    cmpData_length => class_at_0004_cmpData_length,
    mat00_in => class_at_0004_mat00_in,
    mat00_we => class_at_0004_mat00_we,
    mat00_out => class_at_0004_mat00_out,
    mat01_in => class_at_0004_mat01_in,
    mat01_we => class_at_0004_mat01_we,
    mat01_out => class_at_0004_mat01_out,
    mat02_in => class_at_0004_mat02_in,
    mat02_we => class_at_0004_mat02_we,
    mat02_out => class_at_0004_mat02_out,
    mat10_in => class_at_0004_mat10_in,
    mat10_we => class_at_0004_mat10_we,
    mat10_out => class_at_0004_mat10_out,
    mat11_in => class_at_0004_mat11_in,
    mat11_we => class_at_0004_mat11_we,
    mat11_out => class_at_0004_mat11_out,
    mat12_in => class_at_0004_mat12_in,
    mat12_we => class_at_0004_mat12_we,
    mat12_out => class_at_0004_mat12_out,
    modeInterpolation_in => class_at_0004_modeInterpolation_in,
    modeInterpolation_we => class_at_0004_modeInterpolation_we,
    modeInterpolation_out => class_at_0004_modeInterpolation_out,
    modeCompare_in => class_at_0004_modeCompare_in,
    modeCompare_we => class_at_0004_modeCompare_we,
    modeCompare_out => class_at_0004_modeCompare_out,
    diffCompare_in => class_at_0004_diffCompare_in,
    diffCompare_we => class_at_0004_diffCompare_we,
    diffCompare_out => class_at_0004_diffCompare_out,
    clear_busy => class_at_0004_clear_busy,
    clear_req => class_at_0004_clear_req,
    proc_busy => class_at_0004_proc_busy,
    proc_req => class_at_0004_proc_req
  );


end RTL;
